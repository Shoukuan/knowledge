* Path and file = D:\Work\02_SIwave\07_CPA_Flow\A025 PCB RLC Extraction\PCB RLC Extraction.siwaveresults\0002_CPA_Sim_3\0002_CPA_Sim_3_PDN_Channel\0002_CPA_Sim_3_C83410-012_C3L17.sp

.subckt a0002_CPA_Sim_3_C83410-012_C3L17
+ 1 2
C1 1 2 1.000000e-06
.ends a0002_CPA_Sim_3_C83410-012_C3L17
