* contains one subcircuit for each unique part in design

.subckt 602433_081 1 2
C1 1 2 2.200000e-05
.ends 602433_081

.subckt A36096_108 1 2
C1 1 2 1.000000e-05
.ends A36096_108

.subckt C83410_012 1 2
C1 1 2 1.000000e-06
.ends C83410_012

.subckt C97875_001 1 2
C1 1 2 2.200000e-05
.ends C97875_001

.subckt E16347_001 1 2
C1 1 2 1.000000e-08
.ends E16347_001

