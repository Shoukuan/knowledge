* Wide band Macro model for project = 0002_CPA_Sim_3

* Remove the _WB from the file name to use it.
* This file is invalid if spiceModel_WT.sp is not present in the same folder

.include spiceModel_WT.sp

.subckt a0002_CPA_Sim_3
+ U2A5_GND_Group Group_602433-081_C2B2_GND_1 Group_602433-081_C3B10_GND_1
+ Group_A36096-108_C3L22_GND_1 Group_C83410-012_C3L15_GND_1
+ Group_C83410-012_C3L17_GND_1 Group_C83410-012_C3L18_GND_1
+ Group_C83410-012_C3L20_GND_1 Group_C83410-012_C3L24_GND_1
+ Group_C83410-012_C3L26_GND_1 Group_C83410-012_C3L28_GND_1
+ Group_C83410-012_C3L29_GND_1 Group_C97875-001_C3B11_GND_1
+ Group_C97875-001_C3B9_GND_1 Group_E16347-001_C2B12_GND_1
+ Group_E16347-001_C3B17_GND_1 U2A5_V1P0_S0_Group Group_602433-081_C2B2_V1P0_S0_2
+ Group_602433-081_C3B10_V1P0_S0_2 Group_A36096-108_C3L22_V1P0_S0_2
+ Group_C83410-012_C3L15_V1P0_S0_2 Group_C83410-012_C3L17_V1P0_S0_2
+ Group_C83410-012_C3L18_V1P0_S0_2 Group_C83410-012_C3L20_V1P0_S0_2
+ Group_C83410-012_C3L24_V1P0_S0_2 Group_C83410-012_C3L26_V1P0_S0_2
+ Group_C83410-012_C3L28_V1P0_S0_2 Group_C83410-012_C3L29_V1P0_S0_2
+ Group_C97875-001_C3B11_V1P0_S0_2 Group_C97875-001_C3B9_V1P0_S0_2
+ Group_E16347-001_C2B12_V1P0_S0_2 Group_E16347-001_C3B17_V1P0_S0_2
+ XW_V1P0_S0_SINK_ XW_GND_SINK_

V0 Group_602433-081_C2B2_GND_1 0 0.0
V1 Group_602433-081_C3B10_GND_1 0 0.0
V2 Group_A36096-108_C3L22_GND_1 0 0.0
V3 Group_C83410-012_C3L15_GND_1 0 0.0
V4 Group_C83410-012_C3L17_GND_1 0 0.0
V5 Group_C83410-012_C3L18_GND_1 0 0.0
V6 Group_C83410-012_C3L20_GND_1 0 0.0
V7 Group_C83410-012_C3L24_GND_1 0 0.0
V8 Group_C83410-012_C3L26_GND_1 0 0.0
V9 Group_C83410-012_C3L28_GND_1 0 0.0
V10 Group_C83410-012_C3L29_GND_1 0 0.0
V11 Group_C97875-001_C3B11_GND_1 0 0.0
V12 Group_C97875-001_C3B9_GND_1 0 0.0
V13 Group_E16347-001_C2B12_GND_1 0 0.0
V14 Group_E16347-001_C3B17_GND_1 0 0.0


xpackage
+ U2A5_GND_Group U2A5_V1P0_S0_Group Group_602433-081_C2B2_V1P0_S0_2
+ Group_602433-081_C3B10_V1P0_S0_2 Group_A36096-108_C3L22_V1P0_S0_2
+ Group_C83410-012_C3L15_V1P0_S0_2 Group_C83410-012_C3L17_V1P0_S0_2
+ Group_C83410-012_C3L18_V1P0_S0_2 Group_C83410-012_C3L20_V1P0_S0_2
+ Group_C83410-012_C3L24_V1P0_S0_2 Group_C83410-012_C3L26_V1P0_S0_2
+ Group_C83410-012_C3L28_V1P0_S0_2 Group_C83410-012_C3L29_V1P0_S0_2
+ Group_C97875-001_C3B11_V1P0_S0_2 Group_C97875-001_C3B9_V1P0_S0_2
+ Group_E16347-001_C2B12_V1P0_S0_2 Group_E16347-001_C3B17_V1P0_S0_2 XW_GND_SINK_
+ XW_V1P0_S0_SINK_
+ package
.ends a0002_CPA_Sim_3
