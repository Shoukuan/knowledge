* contains one subcircuit for each unique part in design

.subckt G98327_001 1 2
R1 1 2 3.240000e+01
.ends G98327_001

.subckt 602433_081 1 2
C1 1 2 2.200000e-05
.ends 602433_081

.subckt A93548_034 1 2
R1 1 2 1.000000e+04
.ends A93548_034

.subckt A93548_127 1 2
R1 1 2 1.580000e+05
.ends A93548_127

.subckt A36096_108 1 2
C1 1 2 1.000000e-05
.ends A36096_108

.subckt C83410_012 1 2
C1 1 2 1.000000e-06
.ends C83410_012

.subckt A36096_046 1 2
C1 1 2 1.000000e-09
.ends A36096_046

.subckt A36094_025 1 2
C1 1 2 1.000000e-11
.ends A36094_025

.subckt 602433_026 1 2
C1 1 2 2.200000e-06
.ends 602433_026

.subckt A36096_066 1 2
C1 1 2 4.700000e-09
.ends A36096_066

.subckt A93548_056 1 2
R1 1 2 2.260000e+01
.ends A93548_056

.subckt A93548_224 1 2
R1 1 2 4.530000e+04
.ends A93548_224

.subckt E78606_001 1 2
R1 1 2 8.060000e+03
.ends E78606_001

.subckt 602433_075 1 2
C1 1 2 1.000000e-05
.ends 602433_075

.subckt A93548_479 1 2
R1 1 2 1.800000e+05
.ends A93548_479

.subckt G85288_001 1 2
R1 1 2 3.400000e+01
.ends G85288_001

.subckt C97875_001 1 2
C1 1 2 2.200000e-05
.ends C97875_001

.subckt A93548_014 1 2
R1 1 2 1.500000e+03
.ends A93548_014

.subckt 644066_115 1 2
C1 1 2 4.700000e-05
.ends 644066_115

.subckt E57936_001 1 2
C1 1 2 1.000000e-05
.ends E57936_001

.subckt A93548_339 1 2
R1 1 2 1.270000e+04
.ends A93548_339

.subckt A93548_433 1 2
R1 1 2 1.470000e+05
.ends A93548_433

.subckt A93548_248 1 2
R1 1 2 2.740000e+02
.ends A93548_248

.subckt A93548_045 1 2
R1 1 2 4.990000e+01
.ends A93548_045

.subckt A36096_027 1 2
C1 1 2 1.000000e-06
.ends A36096_027

.subckt C17927_001 1 2
R1 1 2 1.000000e-05
.ends C17927_001

.subckt A36095_042 1 2
C1 1 2 1.800000e-11
.ends A36095_042

.subckt A36096_030 1 2
C1 1 2 1.000000e-07
.ends A36096_030

.subckt E16347_001 1 2
C1 1 2 1.000000e-08
.ends E16347_001

.subckt 602433_057 1 2
C1 1 2 4.700000e-08
.ends 602433_057

.subckt A32422_019 1 2
L1 1 2 1.000000e-09
.ends A32422_019

.subckt A93549_023 1 2
R1 1 2 1.000000e+04
.ends A93549_023

.subckt E41735_001 1 2
R1 1 2 4.020000e+04
.ends E41735_001

