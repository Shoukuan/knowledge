* Path and file = D:\Persional\02 SIwave\07 CPA\Workflow\CPA Radhawk RLGC.siwaveresults\0000_CPA_Sim_1\0000_CPA_Sim_1_PDN_Channel\0000_CPA_Sim_1_COMP1_part_COMP1.sp

.subckt a0000_CPA_Sim_1_COMP1_part_COMP1
+ 1 2
C1 1 2 1.000000e-08
.ends a0000_CPA_Sim_1_COMP1_part_COMP1
