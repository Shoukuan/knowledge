* Path and file = D:\Persional\02 SIwave\07 CPA\Workflow\CPA IBIS RLGC.siwaveresults\0000_CPA_Sim_1\0000_CPA_Sim_1_PDN_Channel\0000_CPA_Sim_1_CSP_BGA_BGA.sp

.subckt a0000_CPA_Sim_1_CSP_BGA_BGA
+ BGA_VSS_Group_SINK_ BGA_TXDATA2-_Group_SINK_ BGA_TXDATA2+_Group_SINK_
+ BGA_TXDATA1-_Group_SINK_ BGA_TXDATA5-_Group_SINK_ BGA_TXDATA3+_Group_SINK_
+ BGA_TXDATA7+_Group_SINK_ BGA_TXDATA1+_Group_SINK_ BGA_TXDATA0-_Group_SINK_
+ BGA_TXDATA3-_Group_SINK_ BGA_TXDATA4-_Group_SINK_ BGA_TXDATA4+_Group_SINK_
+ BGA_TXDATA5+_Group_SINK_ BGA_TXDATA6-_Group_SINK_ BGA_TXDATA6+_Group_SINK_
+ BGA_TXDATA7-_Group_SINK_ BGA_RXDATA2+_Group_SINK_ BGA_RXDATA0+_Group_SINK_
+ BGA_RXDATA3+_Group_SINK_ BGA_RXDATA5+_Group_SINK_ BGA_RXDATA1-_Group_SINK_
+ BGA_RXDATA2-_Group_SINK_ BGA_RXDATA0-_Group_SINK_ BGA_RXDATA1+_Group_SINK_
+ BGA_RXDATA3-_Group_SINK_ BGA_RXDATA4+_Group_SINK_ BGA_RXDATA4-_Group_SINK_
+ BGA_RXDATA7+_Group_SINK_ BGA_RXDATA6-_Group_SINK_ BGA_RXDATA5-_Group_SINK_
+ BGA_RXDATA6+_Group_SINK_ BGA_RXDATA7-_Group_SINK_ BGA_TXDATA0+_Group_SINK_
V1 BGA_TXDATA0+_Group_SINK_ 0 1.500000e+00
V2 BGA_RXDATA7-_Group_SINK_ 0 1.500000e+00
V3 BGA_RXDATA6+_Group_SINK_ 0 1.500000e+00
V4 BGA_RXDATA5-_Group_SINK_ 0 1.500000e+00
V5 BGA_RXDATA6-_Group_SINK_ 0 1.500000e+00
V6 BGA_RXDATA7+_Group_SINK_ 0 1.500000e+00
V7 BGA_RXDATA4-_Group_SINK_ 0 1.500000e+00
V8 BGA_RXDATA4+_Group_SINK_ 0 1.500000e+00
V9 BGA_RXDATA3-_Group_SINK_ 0 1.500000e+00
V10 BGA_RXDATA1+_Group_SINK_ 0 1.500000e+00
V11 BGA_RXDATA0-_Group_SINK_ 0 1.500000e+00
V12 BGA_RXDATA2-_Group_SINK_ 0 1.500000e+00
V13 BGA_RXDATA1-_Group_SINK_ 0 1.500000e+00
V14 BGA_RXDATA5+_Group_SINK_ 0 1.500000e+00
V15 BGA_RXDATA3+_Group_SINK_ 0 1.500000e+00
V16 BGA_RXDATA0+_Group_SINK_ 0 1.500000e+00
V17 BGA_RXDATA2+_Group_SINK_ 0 1.500000e+00
V18 BGA_TXDATA7-_Group_SINK_ 0 1.500000e+00
V19 BGA_TXDATA6+_Group_SINK_ 0 1.500000e+00
V20 BGA_TXDATA6-_Group_SINK_ 0 1.500000e+00
V21 BGA_TXDATA5+_Group_SINK_ 0 1.500000e+00
V22 BGA_TXDATA4+_Group_SINK_ 0 1.500000e+00
V23 BGA_TXDATA4-_Group_SINK_ 0 1.500000e+00
V24 BGA_TXDATA3-_Group_SINK_ 0 1.500000e+00
V25 BGA_TXDATA0-_Group_SINK_ 0 1.500000e+00
V26 BGA_TXDATA1+_Group_SINK_ 0 1.500000e+00
V27 BGA_TXDATA7+_Group_SINK_ 0 1.500000e+00
V28 BGA_TXDATA3+_Group_SINK_ 0 1.500000e+00
V29 BGA_TXDATA5-_Group_SINK_ 0 1.500000e+00
V30 BGA_TXDATA1-_Group_SINK_ 0 1.500000e+00
V31 BGA_TXDATA2+_Group_SINK_ 0 1.500000e+00
V32 BGA_TXDATA2-_Group_SINK_ 0 1.500000e+00
V33 BGA_VSS_Group_SINK_ 0 0.000000e+00
.ends a0000_CPA_Sim_1_CSP_BGA_BGA
