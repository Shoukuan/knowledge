* Macro model for project = 0000_CPA_Sim_1

.subckt a0000_CPA_Sim_1
+ FCHIP_RXDATA0+_Group FCHIP_RXDATA0-_Group FCHIP_RXDATA1+_Group
+ FCHIP_RXDATA1-_Group FCHIP_RXDATA2+_Group FCHIP_RXDATA2-_Group
+ FCHIP_RXDATA3+_Group FCHIP_RXDATA3-_Group FCHIP_RXDATA4+_Group
+ FCHIP_RXDATA4-_Group FCHIP_RXDATA5+_Group FCHIP_RXDATA5-_Group
+ FCHIP_RXDATA6+_Group FCHIP_RXDATA6-_Group FCHIP_RXDATA7+_Group
+ FCHIP_RXDATA7-_Group FCHIP_TXDATA0+_Group FCHIP_TXDATA0-_Group
+ FCHIP_TXDATA1+_Group FCHIP_TXDATA1-_Group FCHIP_TXDATA2+_Group
+ FCHIP_TXDATA2-_Group FCHIP_TXDATA3+_Group FCHIP_TXDATA3-_Group
+ FCHIP_TXDATA4+_Group FCHIP_TXDATA4-_Group FCHIP_TXDATA5+_Group
+ FCHIP_TXDATA5-_Group FCHIP_TXDATA6+_Group FCHIP_TXDATA6-_Group
+ FCHIP_TXDATA7+_Group FCHIP_TXDATA7-_Group FCHIP_VSS_Group
+ BGA_RXDATA0+_Group_SINK_ BGA_VSS_Group_SINK_ BGA_RXDATA0-_Group_SINK_
+ BGA_RXDATA1+_Group_SINK_ BGA_RXDATA1-_Group_SINK_ BGA_RXDATA2+_Group_SINK_
+ BGA_RXDATA2-_Group_SINK_ BGA_RXDATA3+_Group_SINK_ BGA_RXDATA3-_Group_SINK_
+ BGA_RXDATA4+_Group_SINK_ BGA_RXDATA4-_Group_SINK_ BGA_RXDATA5+_Group_SINK_
+ BGA_RXDATA5-_Group_SINK_ BGA_RXDATA6+_Group_SINK_ BGA_RXDATA6-_Group_SINK_
+ BGA_RXDATA7+_Group_SINK_ BGA_RXDATA7-_Group_SINK_ BGA_TXDATA0+_Group_SINK_
+ BGA_TXDATA0-_Group_SINK_ BGA_TXDATA1+_Group_SINK_ BGA_TXDATA1-_Group_SINK_
+ BGA_TXDATA2+_Group_SINK_ BGA_TXDATA2-_Group_SINK_ BGA_TXDATA3+_Group_SINK_
+ BGA_TXDATA3-_Group_SINK_ BGA_TXDATA4+_Group_SINK_ BGA_TXDATA4-_Group_SINK_
+ BGA_TXDATA5+_Group_SINK_ BGA_TXDATA5-_Group_SINK_ BGA_TXDATA6+_Group_SINK_
+ BGA_TXDATA6-_Group_SINK_ BGA_TXDATA7+_Group_SINK_ BGA_TXDATA7-_Group_SINK_

L1_0_0 FCHIP_RXDATA0+_Group FCHIP_RXDATA0+_Group_mid 9.905112e-10
L2_0_0 FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA0+_Group_resist 9.905112e-10
L1_1_1 FCHIP_RXDATA0-_Group FCHIP_RXDATA0-_Group_mid 1.162018e-09
L2_1_1 FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA0-_Group_resist 1.162018e-09
L1_2_2 FCHIP_RXDATA1+_Group FCHIP_RXDATA1+_Group_mid 1.334631e-09
L2_2_2 FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA1+_Group_resist 1.334631e-09
L1_3_3 FCHIP_RXDATA1-_Group FCHIP_RXDATA1-_Group_mid 1.299891e-09
L2_3_3 FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA1-_Group_resist 1.299891e-09
L1_4_4 FCHIP_RXDATA2+_Group FCHIP_RXDATA2+_Group_mid 1.197885e-09
L2_4_4 FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA2+_Group_resist 1.197885e-09
L1_5_5 FCHIP_RXDATA2-_Group FCHIP_RXDATA2-_Group_mid 1.264490e-09
L2_5_5 FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA2-_Group_resist 1.264490e-09
L1_6_6 FCHIP_RXDATA3+_Group FCHIP_RXDATA3+_Group_mid 1.089192e-09
L2_6_6 FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA3+_Group_resist 1.089192e-09
L1_7_7 FCHIP_RXDATA3-_Group FCHIP_RXDATA3-_Group_mid 1.082448e-09
L2_7_7 FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA3-_Group_resist 1.082448e-09
L1_8_8 FCHIP_RXDATA4+_Group FCHIP_RXDATA4+_Group_mid 1.254567e-09
L2_8_8 FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA4+_Group_resist 1.254567e-09
L1_9_9 FCHIP_RXDATA4-_Group FCHIP_RXDATA4-_Group_mid 1.238376e-09
L2_9_9 FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA4-_Group_resist 1.238376e-09
L1_10_10 FCHIP_RXDATA5+_Group FCHIP_RXDATA5+_Group_mid 1.385218e-09
L2_10_10 FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA5+_Group_resist 1.385218e-09
L1_11_11 FCHIP_RXDATA5-_Group FCHIP_RXDATA5-_Group_mid 1.207817e-09
L2_11_11 FCHIP_RXDATA5-_Group_mid FCHIP_RXDATA5-_Group_resist 1.207817e-09
L1_12_12 FCHIP_RXDATA6+_Group FCHIP_RXDATA6+_Group_mid 1.156606e-09
L2_12_12 FCHIP_RXDATA6+_Group_mid FCHIP_RXDATA6+_Group_resist 1.156606e-09
L1_13_13 FCHIP_RXDATA6-_Group FCHIP_RXDATA6-_Group_mid 1.181862e-09
L2_13_13 FCHIP_RXDATA6-_Group_mid FCHIP_RXDATA6-_Group_resist 1.181862e-09
L1_14_14 FCHIP_RXDATA7+_Group FCHIP_RXDATA7+_Group_mid 1.299681e-09
L2_14_14 FCHIP_RXDATA7+_Group_mid FCHIP_RXDATA7+_Group_resist 1.299681e-09
L1_15_15 FCHIP_RXDATA7-_Group FCHIP_RXDATA7-_Group_mid 1.231099e-09
L2_15_15 FCHIP_RXDATA7-_Group_mid FCHIP_RXDATA7-_Group_resist 1.231099e-09
L1_16_16 FCHIP_TXDATA0+_Group FCHIP_TXDATA0+_Group_mid 1.014526e-09
L2_16_16 FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA0+_Group_resist 1.014526e-09
L1_17_17 FCHIP_TXDATA0-_Group FCHIP_TXDATA0-_Group_mid 1.145957e-09
L2_17_17 FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA0-_Group_resist 1.145957e-09
L1_18_18 FCHIP_TXDATA1+_Group FCHIP_TXDATA1+_Group_mid 1.188322e-09
L2_18_18 FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA1+_Group_resist 1.188322e-09
L1_19_19 FCHIP_TXDATA1-_Group FCHIP_TXDATA1-_Group_mid 1.183384e-09
L2_19_19 FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA1-_Group_resist 1.183384e-09
L1_20_20 FCHIP_TXDATA2+_Group FCHIP_TXDATA2+_Group_mid 1.223772e-09
L2_20_20 FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA2+_Group_resist 1.223772e-09
L1_21_21 FCHIP_TXDATA2-_Group FCHIP_TXDATA2-_Group_mid 1.208193e-09
L2_21_21 FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA2-_Group_resist 1.208193e-09
L1_22_22 FCHIP_TXDATA3+_Group FCHIP_TXDATA3+_Group_mid 1.041089e-09
L2_22_22 FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA3+_Group_resist 1.041089e-09
L1_23_23 FCHIP_TXDATA3-_Group FCHIP_TXDATA3-_Group_mid 1.065559e-09
L2_23_23 FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA3-_Group_resist 1.065559e-09
L1_24_24 FCHIP_TXDATA4+_Group FCHIP_TXDATA4+_Group_mid 1.226584e-09
L2_24_24 FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA4+_Group_resist 1.226584e-09
L1_25_25 FCHIP_TXDATA4-_Group FCHIP_TXDATA4-_Group_mid 1.257641e-09
L2_25_25 FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA4-_Group_resist 1.257641e-09
L1_26_26 FCHIP_TXDATA5+_Group FCHIP_TXDATA5+_Group_mid 1.416330e-09
L2_26_26 FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA5+_Group_resist 1.416330e-09
L1_27_27 FCHIP_TXDATA5-_Group FCHIP_TXDATA5-_Group_mid 1.238625e-09
L2_27_27 FCHIP_TXDATA5-_Group_mid FCHIP_TXDATA5-_Group_resist 1.238625e-09
L1_28_28 FCHIP_TXDATA6+_Group FCHIP_TXDATA6+_Group_mid 1.218246e-09
L2_28_28 FCHIP_TXDATA6+_Group_mid FCHIP_TXDATA6+_Group_resist 1.218246e-09
L1_29_29 FCHIP_TXDATA6-_Group FCHIP_TXDATA6-_Group_mid 1.176811e-09
L2_29_29 FCHIP_TXDATA6-_Group_mid FCHIP_TXDATA6-_Group_resist 1.176811e-09
L1_30_30 FCHIP_TXDATA7+_Group FCHIP_TXDATA7+_Group_mid 1.202187e-09
L2_30_30 FCHIP_TXDATA7+_Group_mid FCHIP_TXDATA7+_Group_resist 1.202187e-09
L1_31_31 FCHIP_TXDATA7-_Group FCHIP_TXDATA7-_Group_mid 1.297676e-09
L2_31_31 FCHIP_TXDATA7-_Group_mid FCHIP_TXDATA7-_Group_resist 1.297676e-09
L1_32_32 FCHIP_VSS_Group FCHIP_VSS_Group_mid 5.000000e-17
L2_32_32 FCHIP_VSS_Group_mid FCHIP_VSS_Group_resist 5.000000e-17


R_d_1 FCHIP_RXDATA0+_Group_resist BGA_RXDATA0+_Group_SINK_ 3.770891e-02
R_d_2 FCHIP_RXDATA0-_Group_resist BGA_RXDATA0-_Group_SINK_ 4.001462e-02
R_d_3 FCHIP_RXDATA1+_Group_resist BGA_RXDATA1+_Group_SINK_ 4.219923e-02
R_d_4 FCHIP_RXDATA1-_Group_resist BGA_RXDATA1-_Group_SINK_ 4.022461e-02
R_d_5 FCHIP_RXDATA2+_Group_resist BGA_RXDATA2+_Group_SINK_ 3.590737e-02
R_d_6 FCHIP_RXDATA2-_Group_resist BGA_RXDATA2-_Group_SINK_ 3.662762e-02
R_d_7 FCHIP_RXDATA3+_Group_resist BGA_RXDATA3+_Group_SINK_ 3.275829e-02
R_d_8 FCHIP_RXDATA3-_Group_resist BGA_RXDATA3-_Group_SINK_ 3.326557e-02
R_d_9 FCHIP_RXDATA4+_Group_resist BGA_RXDATA4+_Group_SINK_ 4.033628e-02
R_d_10 FCHIP_RXDATA4-_Group_resist BGA_RXDATA4-_Group_SINK_ 3.978307e-02
R_d_11 FCHIP_RXDATA5+_Group_resist BGA_RXDATA5+_Group_SINK_ 5.098034e-02
R_d_12 FCHIP_RXDATA5-_Group_resist BGA_RXDATA5-_Group_SINK_ 5.065322e-02
R_d_13 FCHIP_RXDATA6+_Group_resist BGA_RXDATA6+_Group_SINK_ 3.001861e-02
R_d_14 FCHIP_RXDATA6-_Group_resist BGA_RXDATA6-_Group_SINK_ 3.103480e-02
R_d_15 FCHIP_RXDATA7+_Group_resist BGA_RXDATA7+_Group_SINK_ 3.566011e-02
R_d_16 FCHIP_RXDATA7-_Group_resist BGA_RXDATA7-_Group_SINK_ 3.317870e-02
R_d_17 FCHIP_TXDATA0+_Group_resist BGA_TXDATA0+_Group_SINK_ 3.746788e-02
R_d_18 FCHIP_TXDATA0-_Group_resist BGA_TXDATA0-_Group_SINK_ 3.972360e-02
R_d_19 FCHIP_TXDATA1+_Group_resist BGA_TXDATA1+_Group_SINK_ 4.067288e-02
R_d_20 FCHIP_TXDATA1-_Group_resist BGA_TXDATA1-_Group_SINK_ 4.203842e-02
R_d_21 FCHIP_TXDATA2+_Group_resist BGA_TXDATA2+_Group_SINK_ 3.965275e-02
R_d_22 FCHIP_TXDATA2-_Group_resist BGA_TXDATA2-_Group_SINK_ 3.927664e-02
R_d_23 FCHIP_TXDATA3+_Group_resist BGA_TXDATA3+_Group_SINK_ 3.325824e-02
R_d_24 FCHIP_TXDATA3-_Group_resist BGA_TXDATA3-_Group_SINK_ 3.300170e-02
R_d_25 FCHIP_TXDATA4+_Group_resist BGA_TXDATA4+_Group_SINK_ 3.867945e-02
R_d_26 FCHIP_TXDATA4-_Group_resist BGA_TXDATA4-_Group_SINK_ 3.892028e-02
R_d_27 FCHIP_TXDATA5+_Group_resist BGA_TXDATA5+_Group_SINK_ 5.114009e-02
R_d_28 FCHIP_TXDATA5-_Group_resist BGA_TXDATA5-_Group_SINK_ 5.092169e-02
R_d_29 FCHIP_TXDATA6+_Group_resist BGA_TXDATA6+_Group_SINK_ 3.104464e-02
R_d_30 FCHIP_TXDATA6-_Group_resist BGA_TXDATA6-_Group_SINK_ 3.054399e-02
R_d_31 FCHIP_TXDATA7+_Group_resist BGA_TXDATA7+_Group_SINK_ 3.223324e-02
R_d_32 FCHIP_TXDATA7-_Group_resist BGA_TXDATA7-_Group_SINK_ 3.544219e-02
R_d_33 FCHIP_VSS_Group_resist BGA_VSS_Group_SINK_ 4.698643e-05
K1_0_1  L1_0_0  L1_1_1  3.577512e-01
K2_0_1  L2_0_0  L2_1_1  3.577512e-01
K1_0_2  L1_0_0  L1_2_2  2.302114e-02
K2_0_2  L2_0_0  L2_2_2  2.302114e-02
K1_0_3  L1_0_0  L1_3_3  2.642403e-02
K2_0_3  L2_0_0  L2_3_3  2.642403e-02
K1_0_4  L1_0_0  L1_4_4  5.080673e-03
K2_0_4  L2_0_0  L2_4_4  5.080673e-03
K1_0_5  L1_0_0  L1_5_5  6.530930e-03
K2_0_5  L2_0_0  L2_5_5  6.530930e-03
K1_0_6  L1_0_0  L1_6_6  1.041336e-03
K2_0_6  L2_0_0  L2_6_6  1.041336e-03
K1_0_7  L1_0_0  L1_7_7  9.295026e-04
K2_0_7  L2_0_0  L2_7_7  9.295026e-04
K1_0_8  L1_0_0  L1_8_8  7.469485e-04
K2_0_8  L2_0_0  L2_8_8  7.469485e-04
K1_0_9  L1_0_0  L1_9_9  7.833216e-04
K2_0_9  L2_0_0  L2_9_9  7.833216e-04
K1_0_10  L1_0_0  L1_10_10  4.845153e-04
K2_0_10  L2_0_0  L2_10_10  4.845153e-04
K1_0_11  L1_0_0  L1_11_11  5.043174e-04
K2_0_11  L2_0_0  L2_11_11  5.043174e-04
K1_0_12  L1_0_0  L1_12_12  6.053444e-04
K2_0_12  L2_0_0  L2_12_12  6.053444e-04
K1_0_13  L1_0_0  L1_13_13  5.952698e-04
K2_0_13  L2_0_0  L2_13_13  5.952698e-04
K1_0_14  L1_0_0  L1_14_14  5.677314e-04
K2_0_14  L2_0_0  L2_14_14  5.677314e-04
K1_0_15  L1_0_0  L1_15_15  5.936215e-04
K2_0_15  L2_0_0  L2_15_15  5.936215e-04
K1_0_16  L1_0_0  L1_16_16  4.498297e-04
K2_0_16  L2_0_0  L2_16_16  4.498297e-04
K1_0_17  L1_0_0  L1_17_17  5.774148e-04
K2_0_17  L2_0_0  L2_17_17  5.774148e-04
K1_0_18  L1_0_0  L1_18_18  5.914021e-04
K2_0_18  L2_0_0  L2_18_18  5.914021e-04
K1_0_19  L1_0_0  L1_19_19  5.961229e-04
K2_0_19  L2_0_0  L2_19_19  5.961229e-04
K1_0_20  L1_0_0  L1_20_20  6.057647e-04
K2_0_20  L2_0_0  L2_20_20  6.057647e-04
K1_0_21  L1_0_0  L1_21_21  5.998353e-04
K2_0_21  L2_0_0  L2_21_21  5.998353e-04
K1_0_22  L1_0_0  L1_22_22  6.616274e-04
K2_0_22  L2_0_0  L2_22_22  6.616274e-04
K1_0_23  L1_0_0  L1_23_23  6.566995e-04
K2_0_23  L2_0_0  L2_23_23  6.566995e-04
K1_0_24  L1_0_0  L1_24_24  5.999326e-04
K2_0_24  L2_0_0  L2_24_24  5.999326e-04
K1_0_25  L1_0_0  L1_25_25  5.966218e-04
K2_0_25  L2_0_0  L2_25_25  5.966218e-04
K1_0_26  L1_0_0  L1_26_26  5.493427e-04
K2_0_26  L2_0_0  L2_26_26  5.493427e-04
K1_0_27  L1_0_0  L1_27_27  5.519497e-04
K2_0_27  L2_0_0  L2_27_27  5.519497e-04
K1_0_28  L1_0_0  L1_28_28  6.013541e-04
K2_0_28  L2_0_0  L2_28_28  6.013541e-04
K1_0_29  L1_0_0  L1_29_29  6.084127e-04
K2_0_29  L2_0_0  L2_29_29  6.084127e-04
K1_0_30  L1_0_0  L1_30_30  5.967954e-04
K2_0_30  L2_0_0  L2_30_30  5.967954e-04
K1_0_31  L1_0_0  L1_31_31  5.829643e-04
K2_0_31  L2_0_0  L2_31_31  5.829643e-04
K1_1_2  L1_1_1  L1_2_2  4.794070e-02
K2_1_2  L2_1_1  L2_2_2  4.794070e-02
K1_1_3  L1_1_1  L1_3_3  3.548271e-02
K2_1_3  L2_1_1  L2_3_3  3.548271e-02
K1_1_4  L1_1_1  L1_4_4  8.475985e-03
K2_1_4  L2_1_1  L2_4_4  8.475985e-03
K1_1_5  L1_1_1  L1_5_5  1.007640e-02
K2_1_5  L2_1_1  L2_5_5  1.007640e-02
K1_1_6  L1_1_1  L1_6_6  1.562136e-03
K2_1_6  L2_1_1  L2_6_6  1.562136e-03
K1_1_7  L1_1_1  L1_7_7  1.544564e-03
K2_1_7  L2_1_1  L2_7_7  1.544564e-03
K1_1_8  L1_1_1  L1_8_8  9.328669e-04
K2_1_8  L2_1_1  L2_8_8  9.328669e-04
K1_1_9  L1_1_1  L1_9_9  1.031532e-03
K2_1_9  L2_1_1  L2_9_9  1.031532e-03
K1_1_10  L1_1_1  L1_10_10  5.889295e-04
K2_1_10  L2_1_1  L2_10_10  5.889295e-04
K1_1_11  L1_1_1  L1_11_11  6.163218e-04
K2_1_11  L2_1_1  L2_11_11  6.163218e-04
K1_1_12  L1_1_1  L1_12_12  5.459304e-04
K2_1_12  L2_1_1  L2_12_12  5.459304e-04
K1_1_13  L1_1_1  L1_13_13  5.267376e-04
K2_1_13  L2_1_1  L2_13_13  5.267376e-04
K1_1_14  L1_1_1  L1_14_14  4.820728e-04
K2_1_14  L2_1_1  L2_14_14  4.820728e-04
K1_1_15  L1_1_1  L1_15_15  5.263482e-04
K2_1_15  L2_1_1  L2_15_15  5.263482e-04
K1_1_16  L1_1_1  L1_16_16  6.185214e-04
K2_1_16  L2_1_1  L2_16_16  6.185214e-04
K1_1_17  L1_1_1  L1_17_17  5.107314e-04
K2_1_17  L2_1_1  L2_17_17  5.107314e-04
K1_1_18  L1_1_1  L1_18_18  5.533401e-04
K2_1_18  L2_1_1  L2_18_18  5.533401e-04
K1_1_19  L1_1_1  L1_19_19  5.478718e-04
K2_1_19  L2_1_1  L2_19_19  5.478718e-04
K1_1_20  L1_1_1  L1_20_20  5.475471e-04
K2_1_20  L2_1_1  L2_20_20  5.475471e-04
K1_1_21  L1_1_1  L1_21_21  5.507921e-04
K2_1_21  L2_1_1  L2_21_21  5.507921e-04
K1_1_22  L1_1_1  L1_22_22  5.966731e-04
K2_1_22  L2_1_1  L2_22_22  5.966731e-04
K1_1_23  L1_1_1  L1_23_23  5.839342e-04
K2_1_23  L2_1_1  L2_23_23  5.839342e-04
K1_1_24  L1_1_1  L1_24_24  5.395597e-04
K2_1_24  L2_1_1  L2_24_24  5.395597e-04
K1_1_25  L1_1_1  L1_25_25  5.405872e-04
K2_1_25  L2_1_1  L2_25_25  5.405872e-04
K1_1_26  L1_1_1  L1_26_26  5.072601e-04
K2_1_26  L2_1_1  L2_26_26  5.072601e-04
K1_1_27  L1_1_1  L1_27_27  5.195215e-04
K2_1_27  L2_1_1  L2_27_27  5.195215e-04
K1_1_28  L1_1_1  L1_28_28  5.399358e-04
K2_1_28  L2_1_1  L2_28_28  5.399358e-04
K1_1_29  L1_1_1  L1_29_29  5.433627e-04
K2_1_29  L2_1_1  L2_29_29  5.433627e-04
K1_1_30  L1_1_1  L1_30_30  5.301328e-04
K2_1_30  L2_1_1  L2_30_30  5.301328e-04
K1_1_31  L1_1_1  L1_31_31  4.999797e-04
K2_1_31  L2_1_1  L2_31_31  4.999797e-04
K1_2_3  L1_2_2  L1_3_3  4.366806e-01
K2_2_3  L2_2_2  L2_3_3  4.366806e-01
K1_2_4  L1_2_2  L1_4_4  8.208023e-02
K2_2_4  L2_2_2  L2_4_4  8.208023e-02
K1_2_5  L1_2_2  L1_5_5  1.139976e-01
K2_2_5  L2_2_2  L2_5_5  1.139976e-01
K1_2_6  L1_2_2  L1_6_6  1.036941e-02
K2_2_6  L2_2_2  L2_6_6  1.036941e-02
K1_2_7  L1_2_2  L1_7_7  1.165173e-02
K2_2_7  L2_2_2  L2_7_7  1.165173e-02
K1_2_8  L1_2_2  L1_8_8  3.373820e-03
K2_2_8  L2_2_2  L2_8_8  3.373820e-03
K1_2_9  L1_2_2  L1_9_9  4.534554e-03
K2_2_9  L2_2_2  L2_9_9  4.534554e-03
K1_2_10  L1_2_2  L1_10_10  1.523907e-03
K2_2_10  L2_2_2  L2_10_10  1.523907e-03
K1_2_11  L1_2_2  L1_11_11  1.214184e-03
K2_2_11  L2_2_2  L2_11_11  1.214184e-03
K1_2_12  L1_2_2  L1_12_12  6.295708e-04
K2_2_12  L2_2_2  L2_12_12  6.295708e-04
K1_2_13  L1_2_2  L1_13_13  5.755114e-04
K2_2_13  L2_2_2  L2_13_13  5.755114e-04
K1_2_14  L1_2_2  L1_14_14  4.933902e-04
K2_2_14  L2_2_2  L2_14_14  4.933902e-04
K1_2_15  L1_2_2  L1_15_15  5.325008e-04
K2_2_15  L2_2_2  L2_15_15  5.325008e-04
K1_2_16  L1_2_2  L1_16_16  5.609978e-04
K2_2_16  L2_2_2  L2_16_16  5.609978e-04
K1_2_17  L1_2_2  L1_17_17  5.081654e-04
K2_2_17  L2_2_2  L2_17_17  5.081654e-04
K1_2_18  L1_2_2  L1_18_18  5.514374e-04
K2_2_18  L2_2_2  L2_18_18  5.514374e-04
K1_2_19  L1_2_2  L1_19_19  5.432530e-04
K2_2_19  L2_2_2  L2_19_19  5.432530e-04
K1_2_20  L1_2_2  L1_20_20  5.475919e-04
K2_2_20  L2_2_2  L2_20_20  5.475919e-04
K1_2_21  L1_2_2  L1_21_21  5.590087e-04
K2_2_21  L2_2_2  L2_21_21  5.590087e-04
K1_2_22  L1_2_2  L1_22_22  6.058337e-04
K2_2_22  L2_2_2  L2_22_22  6.058337e-04
K1_2_23  L1_2_2  L1_23_23  5.942482e-04
K2_2_23  L2_2_2  L2_23_23  5.942482e-04
K1_2_24  L1_2_2  L1_24_24  5.501591e-04
K2_2_24  L2_2_2  L2_24_24  5.501591e-04
K1_2_25  L1_2_2  L1_25_25  5.422106e-04
K2_2_25  L2_2_2  L2_25_25  5.422106e-04
K1_2_26  L1_2_2  L1_26_26  5.043624e-04
K2_2_26  L2_2_2  L2_26_26  5.043624e-04
K1_2_27  L1_2_2  L1_27_27  5.126920e-04
K2_2_27  L2_2_2  L2_27_27  5.126920e-04
K1_2_28  L1_2_2  L1_28_28  5.384015e-04
K2_2_28  L2_2_2  L2_28_28  5.384015e-04
K1_2_29  L1_2_2  L1_29_29  5.411100e-04
K2_2_29  L2_2_2  L2_29_29  5.411100e-04
K1_2_30  L1_2_2  L1_30_30  5.228482e-04
K2_2_30  L2_2_2  L2_30_30  5.228482e-04
K1_2_31  L1_2_2  L1_31_31  4.923541e-04
K2_2_31  L2_2_2  L2_31_31  4.923541e-04
K1_3_4  L1_3_3  L1_4_4  5.939504e-02
K2_3_4  L2_3_3  L2_4_4  5.939504e-02
K1_3_5  L1_3_3  L1_5_5  8.139549e-02
K2_3_5  L2_3_3  L2_5_5  8.139549e-02
K1_3_6  L1_3_3  L1_6_6  7.304268e-03
K2_3_6  L2_3_3  L2_6_6  7.304268e-03
K1_3_7  L1_3_3  L1_7_7  8.389242e-03
K2_3_7  L2_3_3  L2_7_7  8.389242e-03
K1_3_8  L1_3_3  L1_8_8  2.393615e-03
K2_3_8  L2_3_3  L2_8_8  2.393615e-03
K1_3_9  L1_3_3  L1_9_9  3.067687e-03
K2_3_9  L2_3_3  L2_9_9  3.067687e-03
K1_3_10  L1_3_3  L1_10_10  1.147567e-03
K2_3_10  L2_3_3  L2_10_10  1.147567e-03
K1_3_11  L1_3_3  L1_11_11  9.604216e-04
K2_3_11  L2_3_3  L2_11_11  9.604216e-04
K1_3_12  L1_3_3  L1_12_12  5.975747e-04
K2_3_12  L2_3_3  L2_12_12  5.975747e-04
K1_3_13  L1_3_3  L1_13_13  5.616600e-04
K2_3_13  L2_3_3  L2_13_13  5.616600e-04
K1_3_14  L1_3_3  L1_14_14  5.112560e-04
K2_3_14  L2_3_3  L2_14_14  5.112560e-04
K1_3_15  L1_3_3  L1_15_15  5.236397e-04
K2_3_15  L2_3_3  L2_15_15  5.236397e-04
K1_3_16  L1_3_3  L1_16_16  5.730486e-04
K2_3_16  L2_3_3  L2_16_16  5.730486e-04
K1_3_17  L1_3_3  L1_17_17  5.071474e-04
K2_3_17  L2_3_3  L2_17_17  5.071474e-04
K1_3_18  L1_3_3  L1_18_18  5.557208e-04
K2_3_18  L2_3_3  L2_18_18  5.557208e-04
K1_3_19  L1_3_3  L1_19_19  5.410786e-04
K2_3_19  L2_3_3  L2_19_19  5.410786e-04
K1_3_20  L1_3_3  L1_20_20  5.465769e-04
K2_3_20  L2_3_3  L2_20_20  5.465769e-04
K1_3_21  L1_3_3  L1_21_21  5.572333e-04
K2_3_21  L2_3_3  L2_21_21  5.572333e-04
K1_3_22  L1_3_3  L1_22_22  6.076987e-04
K2_3_22  L2_3_3  L2_22_22  6.076987e-04
K1_3_23  L1_3_3  L1_23_23  5.995732e-04
K2_3_23  L2_3_3  L2_23_23  5.995732e-04
K1_3_24  L1_3_3  L1_24_24  5.546253e-04
K2_3_24  L2_3_3  L2_24_24  5.546253e-04
K1_3_25  L1_3_3  L1_25_25  5.483716e-04
K2_3_25  L2_3_3  L2_25_25  5.483716e-04
K1_3_26  L1_3_3  L1_26_26  5.035145e-04
K2_3_26  L2_3_3  L2_26_26  5.035145e-04
K1_3_27  L1_3_3  L1_27_27  5.082485e-04
K2_3_27  L2_3_3  L2_27_27  5.082485e-04
K1_3_28  L1_3_3  L1_28_28  5.425927e-04
K2_3_28  L2_3_3  L2_28_28  5.425927e-04
K1_3_29  L1_3_3  L1_29_29  5.429466e-04
K2_3_29  L2_3_3  L2_29_29  5.429466e-04
K1_3_30  L1_3_3  L1_30_30  5.293973e-04
K2_3_30  L2_3_3  L2_30_30  5.293973e-04
K1_3_31  L1_3_3  L1_31_31  5.032598e-04
K2_3_31  L2_3_3  L2_31_31  5.032598e-04
K1_4_5  L1_4_4  L1_5_5  4.607233e-01
K2_4_5  L2_4_4  L2_5_5  4.607233e-01
K1_4_6  L1_4_4  L1_6_6  8.396967e-02
K2_4_6  L2_4_4  L2_6_6  8.396967e-02
K1_4_7  L1_4_4  L1_7_7  1.107419e-01
K2_4_7  L2_4_4  L2_7_7  1.107419e-01
K1_4_8  L1_4_4  L1_8_8  1.646741e-02
K2_4_8  L2_4_4  L2_8_8  1.646741e-02
K1_4_9  L1_4_4  L1_9_9  2.354359e-02
K2_4_9  L2_4_4  L2_9_9  2.354359e-02
K1_4_10  L1_4_4  L1_10_10  7.720131e-03
K2_4_10  L2_4_4  L2_10_10  7.720131e-03
K1_4_11  L1_4_4  L1_11_11  4.889340e-03
K2_4_11  L2_4_4  L2_11_11  4.889340e-03
K1_4_12  L1_4_4  L1_12_12  1.344902e-03
K2_4_12  L2_4_4  L2_12_12  1.344902e-03
K1_4_13  L1_4_4  L1_13_13  1.160629e-03
K2_4_13  L2_4_4  L2_13_13  1.160629e-03
K1_4_14  L1_4_4  L1_14_14  7.756281e-04
K2_4_14  L2_4_4  L2_14_14  7.756281e-04
K1_4_15  L1_4_4  L1_15_15  6.821748e-04
K2_4_15  L2_4_4  L2_15_15  6.821748e-04
K1_4_16  L1_4_4  L1_16_16  6.045880e-04
K2_4_16  L2_4_4  L2_16_16  6.045880e-04
K1_4_17  L1_4_4  L1_17_17  5.321572e-04
K2_4_17  L2_4_4  L2_17_17  5.321572e-04
K1_4_18  L1_4_4  L1_18_18  5.764163e-04
K2_4_18  L2_4_4  L2_18_18  5.764163e-04
K1_4_19  L1_4_4  L1_19_19  5.721677e-04
K2_4_19  L2_4_4  L2_19_19  5.721677e-04
K1_4_20  L1_4_4  L1_20_20  5.734954e-04
K2_4_20  L2_4_4  L2_20_20  5.734954e-04
K1_4_21  L1_4_4  L1_21_21  5.806291e-04
K2_4_21  L2_4_4  L2_21_21  5.806291e-04
K1_4_22  L1_4_4  L1_22_22  6.339598e-04
K2_4_22  L2_4_4  L2_22_22  6.339598e-04
K1_4_23  L1_4_4  L1_23_23  6.260440e-04
K2_4_23  L2_4_4  L2_23_23  6.260440e-04
K1_4_24  L1_4_4  L1_24_24  5.800917e-04
K2_4_24  L2_4_4  L2_24_24  5.800917e-04
K1_4_25  L1_4_4  L1_25_25  5.750116e-04
K2_4_25  L2_4_4  L2_25_25  5.750116e-04
K1_4_26  L1_4_4  L1_26_26  5.261681e-04
K2_4_26  L2_4_4  L2_26_26  5.261681e-04
K1_4_27  L1_4_4  L1_27_27  5.344140e-04
K2_4_27  L2_4_4  L2_27_27  5.344140e-04
K1_4_28  L1_4_4  L1_28_28  5.650568e-04
K2_4_28  L2_4_4  L2_28_28  5.650568e-04
K1_4_29  L1_4_4  L1_29_29  5.671483e-04
K2_4_29  L2_4_4  L2_29_29  5.671483e-04
K1_4_30  L1_4_4  L1_30_30  5.539939e-04
K2_4_30  L2_4_4  L2_30_30  5.539939e-04
K1_4_31  L1_4_4  L1_31_31  5.172812e-04
K2_4_31  L2_4_4  L2_31_31  5.172812e-04
K1_5_6  L1_5_5  L1_6_6  6.327429e-02
K2_5_6  L2_5_5  L2_6_6  6.327429e-02
K1_5_7  L1_5_5  L1_7_7  7.936492e-02
K2_5_7  L2_5_5  L2_7_7  7.936492e-02
K1_5_8  L1_5_5  L1_8_8  1.401397e-02
K2_5_8  L2_5_5  L2_8_8  1.401397e-02
K1_5_9  L1_5_5  L1_9_9  1.968906e-02
K2_5_9  L2_5_5  L2_9_9  1.968906e-02
K1_5_10  L1_5_5  L1_10_10  6.182412e-03
K2_5_10  L2_5_5  L2_10_10  6.182412e-03
K1_5_11  L1_5_5  L1_11_11  4.097605e-03
K2_5_11  L2_5_5  L2_11_11  4.097605e-03
K1_5_12  L1_5_5  L1_12_12  1.157227e-03
K2_5_12  L2_5_5  L2_12_12  1.157227e-03
K1_5_13  L1_5_5  L1_13_13  9.672513e-04
K2_5_13  L2_5_5  L2_13_13  9.672513e-04
K1_5_14  L1_5_5  L1_14_14  6.750727e-04
K2_5_14  L2_5_5  L2_14_14  6.750727e-04
K1_5_15  L1_5_5  L1_15_15  6.297220e-04
K2_5_15  L2_5_5  L2_15_15  6.297220e-04
K1_5_16  L1_5_5  L1_16_16  5.786571e-04
K2_5_16  L2_5_5  L2_16_16  5.786571e-04
K1_5_17  L1_5_5  L1_17_17  5.172132e-04
K2_5_17  L2_5_5  L2_17_17  5.172132e-04
K1_5_18  L1_5_5  L1_18_18  5.658384e-04
K2_5_18  L2_5_5  L2_18_18  5.658384e-04
K1_5_19  L1_5_5  L1_19_19  5.547253e-04
K2_5_19  L2_5_5  L2_19_19  5.547253e-04
K1_5_20  L1_5_5  L1_20_20  5.593158e-04
K2_5_20  L2_5_5  L2_20_20  5.593158e-04
K1_5_21  L1_5_5  L1_21_21  5.730372e-04
K2_5_21  L2_5_5  L2_21_21  5.730372e-04
K1_5_22  L1_5_5  L1_22_22  6.237816e-04
K2_5_22  L2_5_5  L2_22_22  6.237816e-04
K1_5_23  L1_5_5  L1_23_23  6.154590e-04
K2_5_23  L2_5_5  L2_23_23  6.154590e-04
K1_5_24  L1_5_5  L1_24_24  5.717019e-04
K2_5_24  L2_5_5  L2_24_24  5.717019e-04
K1_5_25  L1_5_5  L1_25_25  5.594062e-04
K2_5_25  L2_5_5  L2_25_25  5.594062e-04
K1_5_26  L1_5_5  L1_26_26  5.175979e-04
K2_5_26  L2_5_5  L2_26_26  5.175979e-04
K1_5_27  L1_5_5  L1_27_27  5.252297e-04
K2_5_27  L2_5_5  L2_27_27  5.252297e-04
K1_5_28  L1_5_5  L1_28_28  5.535932e-04
K2_5_28  L2_5_5  L2_28_28  5.535932e-04
K1_5_29  L1_5_5  L1_29_29  5.564827e-04
K2_5_29  L2_5_5  L2_29_29  5.564827e-04
K1_5_30  L1_5_5  L1_30_30  5.406642e-04
K2_5_30  L2_5_5  L2_30_30  5.406642e-04
K1_5_31  L1_5_5  L1_31_31  5.113324e-04
K2_5_31  L2_5_5  L2_31_31  5.113324e-04
K1_6_7  L1_6_6  L1_7_7  4.321509e-01
K2_6_7  L2_6_6  L2_7_7  4.321509e-01
K1_6_8  L1_6_6  L1_8_8  9.556248e-02
K2_6_8  L2_6_6  L2_8_8  9.556248e-02
K1_6_9  L1_6_6  L1_9_9  1.416311e-01
K2_6_9  L2_6_6  L2_9_9  1.416311e-01
K1_6_10  L1_6_6  L1_10_10  2.584281e-02
K2_6_10  L2_6_6  L2_10_10  2.584281e-02
K1_6_11  L1_6_6  L1_11_11  1.709333e-02
K2_6_11  L2_6_6  L2_11_11  1.709333e-02
K1_6_12  L1_6_6  L1_12_12  3.346633e-03
K2_6_12  L2_6_6  L2_12_12  3.346633e-03
K1_6_13  L1_6_6  L1_13_13  2.333828e-03
K2_6_13  L2_6_6  L2_13_13  2.333828e-03
K1_6_14  L1_6_6  L1_14_14  1.174561e-03
K2_6_14  L2_6_6  L2_14_14  1.174561e-03
K1_6_15  L1_6_6  L1_15_15  9.863679e-04
K2_6_15  L2_6_6  L2_15_15  9.863679e-04
K1_6_16  L1_6_6  L1_16_16  6.330692e-04
K2_6_16  L2_6_6  L2_16_16  6.330692e-04
K1_6_17  L1_6_6  L1_17_17  5.557745e-04
K2_6_17  L2_6_6  L2_17_17  5.557745e-04
K1_6_18  L1_6_6  L1_18_18  6.063034e-04
K2_6_18  L2_6_6  L2_18_18  6.063034e-04
K1_6_19  L1_6_6  L1_19_19  5.966769e-04
K2_6_19  L2_6_6  L2_19_19  5.966769e-04
K1_6_20  L1_6_6  L1_20_20  6.025478e-04
K2_6_20  L2_6_6  L2_20_20  6.025478e-04
K1_6_21  L1_6_6  L1_21_21  6.166819e-04
K2_6_21  L2_6_6  L2_21_21  6.166819e-04
K1_6_22  L1_6_6  L1_22_22  6.674708e-04
K2_6_22  L2_6_6  L2_22_22  6.674708e-04
K1_6_23  L1_6_6  L1_23_23  6.557447e-04
K2_6_23  L2_6_6  L2_23_23  6.557447e-04
K1_6_24  L1_6_6  L1_24_24  6.081328e-04
K2_6_24  L2_6_6  L2_24_24  6.081328e-04
K1_6_25  L1_6_6  L1_25_25  5.999799e-04
K2_6_25  L2_6_6  L2_25_25  5.999799e-04
K1_6_26  L1_6_6  L1_26_26  5.536977e-04
K2_6_26  L2_6_6  L2_26_26  5.536977e-04
K1_6_27  L1_6_6  L1_27_27  5.567802e-04
K2_6_27  L2_6_6  L2_27_27  5.567802e-04
K1_6_28  L1_6_6  L1_28_28  5.951582e-04
K2_6_28  L2_6_6  L2_28_28  5.951582e-04
K1_6_29  L1_6_6  L1_29_29  5.951562e-04
K2_6_29  L2_6_6  L2_29_29  5.951562e-04
K1_6_30  L1_6_6  L1_30_30  5.809391e-04
K2_6_30  L2_6_6  L2_30_30  5.809391e-04
K1_6_31  L1_6_6  L1_31_31  5.511695e-04
K2_6_31  L2_6_6  L2_31_31  5.511695e-04
K1_7_8  L1_7_7  L1_8_8  7.609195e-02
K2_7_8  L2_7_7  L2_8_8  7.609195e-02
K1_7_9  L1_7_7  L1_9_9  9.930957e-02
K2_7_9  L2_7_7  L2_9_9  9.930957e-02
K1_7_10  L1_7_7  L1_10_10  1.908735e-02
K2_7_10  L2_7_7  L2_10_10  1.908735e-02
K1_7_11  L1_7_7  L1_11_11  1.334436e-02
K2_7_11  L2_7_7  L2_11_11  1.334436e-02
K1_7_12  L1_7_7  L1_12_12  2.547678e-03
K2_7_12  L2_7_7  L2_12_12  2.547678e-03
K1_7_13  L1_7_7  L1_13_13  1.707765e-03
K2_7_13  L2_7_7  L2_13_13  1.707765e-03
K1_7_14  L1_7_7  L1_14_14  9.004635e-04
K2_7_14  L2_7_7  L2_14_14  9.004635e-04
K1_7_15  L1_7_7  L1_15_15  8.528991e-04
K2_7_15  L2_7_7  L2_15_15  8.528991e-04
K1_7_16  L1_7_7  L1_16_16  6.364618e-04
K2_7_16  L2_7_7  L2_16_16  6.364618e-04
K1_7_17  L1_7_7  L1_17_17  5.576996e-04
K2_7_17  L2_7_7  L2_17_17  5.576996e-04
K1_7_18  L1_7_7  L1_18_18  6.080188e-04
K2_7_18  L2_7_7  L2_18_18  6.080188e-04
K1_7_19  L1_7_7  L1_19_19  6.005043e-04
K2_7_19  L2_7_7  L2_19_19  6.005043e-04
K1_7_20  L1_7_7  L1_20_20  6.041032e-04
K2_7_20  L2_7_7  L2_20_20  6.041032e-04
K1_7_21  L1_7_7  L1_21_21  6.142015e-04
K2_7_21  L2_7_7  L2_21_21  6.142015e-04
K1_7_22  L1_7_7  L1_22_22  6.671909e-04
K2_7_22  L2_7_7  L2_22_22  6.671909e-04
K1_7_23  L1_7_7  L1_23_23  6.565844e-04
K2_7_23  L2_7_7  L2_23_23  6.565844e-04
K1_7_24  L1_7_7  L1_24_24  6.080161e-04
K2_7_24  L2_7_7  L2_24_24  6.080161e-04
K1_7_25  L1_7_7  L1_25_25  6.022650e-04
K2_7_25  L2_7_7  L2_25_25  6.022650e-04
K1_7_26  L1_7_7  L1_26_26  5.528508e-04
K2_7_26  L2_7_7  L2_26_26  5.528508e-04
K1_7_27  L1_7_7  L1_27_27  5.582756e-04
K2_7_27  L2_7_7  L2_27_27  5.582756e-04
K1_7_28  L1_7_7  L1_28_28  5.952572e-04
K2_7_28  L2_7_7  L2_28_28  5.952572e-04
K1_7_29  L1_7_7  L1_29_29  5.961224e-04
K2_7_29  L2_7_7  L2_29_29  5.961224e-04
K1_7_30  L1_7_7  L1_30_30  5.814280e-04
K2_7_30  L2_7_7  L2_30_30  5.814280e-04
K1_7_31  L1_7_7  L1_31_31  5.495077e-04
K2_7_31  L2_7_7  L2_31_31  5.495077e-04
K1_8_9  L1_8_8  L1_9_9  4.278114e-01
K2_8_9  L2_8_8  L2_9_9  4.278114e-01
K1_8_10  L1_8_8  L1_10_10  1.303058e-01
K2_8_10  L2_8_8  L2_10_10  1.303058e-01
K1_8_11  L1_8_8  L1_11_11  7.679043e-02
K2_8_11  L2_8_8  L2_11_11  7.679043e-02
K1_8_12  L1_8_8  L1_12_12  2.354612e-02
K2_8_12  L2_8_8  L2_12_12  2.354612e-02
K1_8_13  L1_8_8  L1_13_13  1.447400e-02
K2_8_13  L2_8_8  L2_13_13  1.447400e-02
K1_8_14  L1_8_8  L1_14_14  5.507947e-03
K2_8_14  L2_8_8  L2_14_14  5.507947e-03
K1_8_15  L1_8_8  L1_15_15  3.697196e-03
K2_8_15  L2_8_8  L2_15_15  3.697196e-03
K1_8_16  L1_8_8  L1_16_16  5.857268e-04
K2_8_16  L2_8_8  L2_16_16  5.857268e-04
K1_8_17  L1_8_8  L1_17_17  5.152213e-04
K2_8_17  L2_8_8  L2_17_17  5.152213e-04
K1_8_18  L1_8_8  L1_18_18  5.581211e-04
K2_8_18  L2_8_8  L2_18_18  5.581211e-04
K1_8_19  L1_8_8  L1_19_19  5.526619e-04
K2_8_19  L2_8_8  L2_19_19  5.526619e-04
K1_8_20  L1_8_8  L1_20_20  5.577392e-04
K2_8_20  L2_8_8  L2_20_20  5.577392e-04
K1_8_21  L1_8_8  L1_21_21  5.689950e-04
K2_8_21  L2_8_8  L2_21_21  5.689950e-04
K1_8_22  L1_8_8  L1_22_22  6.175180e-04
K2_8_22  L2_8_8  L2_22_22  6.175180e-04
K1_8_23  L1_8_8  L1_23_23  6.081326e-04
K2_8_23  L2_8_8  L2_23_23  6.081326e-04
K1_8_24  L1_8_8  L1_24_24  5.647217e-04
K2_8_24  L2_8_8  L2_24_24  5.647217e-04
K1_8_25  L1_8_8  L1_25_25  5.551051e-04
K2_8_25  L2_8_8  L2_25_25  5.551051e-04
K1_8_26  L1_8_8  L1_26_26  5.139124e-04
K2_8_26  L2_8_8  L2_26_26  5.139124e-04
K1_8_27  L1_8_8  L1_27_27  5.166535e-04
K2_8_27  L2_8_8  L2_27_27  5.166535e-04
K1_8_28  L1_8_8  L1_28_28  5.529432e-04
K2_8_28  L2_8_8  L2_28_28  5.529432e-04
K1_8_29  L1_8_8  L1_29_29  5.539057e-04
K2_8_29  L2_8_8  L2_29_29  5.539057e-04
K1_8_30  L1_8_8  L1_30_30  5.423130e-04
K2_8_30  L2_8_8  L2_30_30  5.423130e-04
K1_8_31  L1_8_8  L1_31_31  5.151594e-04
K2_8_31  L2_8_8  L2_31_31  5.151594e-04
K1_9_10  L1_9_9  L1_10_10  9.158689e-02
K2_9_10  L2_9_9  L2_10_10  9.158689e-02
K1_9_11  L1_9_9  L1_11_11  5.671534e-02
K2_9_11  L2_9_9  L2_11_11  5.671534e-02
K1_9_12  L1_9_9  L1_12_12  1.707424e-02
K2_9_12  L2_9_9  L2_12_12  1.707424e-02
K1_9_13  L1_9_9  L1_13_13  1.005690e-02
K2_9_13  L2_9_9  L2_13_13  1.005690e-02
K1_9_14  L1_9_9  L1_14_14  3.631393e-03
K2_9_14  L2_9_9  L2_14_14  3.631393e-03
K1_9_15  L1_9_9  L1_15_15  2.726782e-03
K2_9_15  L2_9_9  L2_15_15  2.726782e-03
K1_9_16  L1_9_9  L1_16_16  5.848076e-04
K2_9_16  L2_9_9  L2_16_16  5.848076e-04
K1_9_17  L1_9_9  L1_17_17  5.208427e-04
K2_9_17  L2_9_9  L2_17_17  5.208427e-04
K1_9_18  L1_9_9  L1_18_18  5.618793e-04
K2_9_18  L2_9_9  L2_18_18  5.618793e-04
K1_9_19  L1_9_9  L1_19_19  5.569420e-04
K2_9_19  L2_9_9  L2_19_19  5.569420e-04
K1_9_20  L1_9_9  L1_20_20  5.611360e-04
K2_9_20  L2_9_9  L2_20_20  5.611360e-04
K1_9_21  L1_9_9  L1_21_21  5.739041e-04
K2_9_21  L2_9_9  L2_21_21  5.739041e-04
K1_9_22  L1_9_9  L1_22_22  6.230742e-04
K2_9_22  L2_9_9  L2_22_22  6.230742e-04
K1_9_23  L1_9_9  L1_23_23  6.143398e-04
K2_9_23  L2_9_9  L2_23_23  6.143398e-04
K1_9_24  L1_9_9  L1_24_24  5.726557e-04
K2_9_24  L2_9_9  L2_24_24  5.726557e-04
K1_9_25  L1_9_9  L1_25_25  5.604078e-04
K2_9_25  L2_9_9  L2_25_25  5.604078e-04
K1_9_26  L1_9_9  L1_26_26  5.207908e-04
K2_9_26  L2_9_9  L2_26_26  5.207908e-04
K1_9_27  L1_9_9  L1_27_27  5.192430e-04
K2_9_27  L2_9_9  L2_27_27  5.192430e-04
K1_9_28  L1_9_9  L1_28_28  5.585010e-04
K2_9_28  L2_9_9  L2_28_28  5.585010e-04
K1_9_29  L1_9_9  L1_29_29  5.570749e-04
K2_9_29  L2_9_9  L2_29_29  5.570749e-04
K1_9_30  L1_9_9  L1_30_30  5.464087e-04
K2_9_30  L2_9_9  L2_30_30  5.464087e-04
K1_9_31  L1_9_9  L1_31_31  5.188803e-04
K2_9_31  L2_9_9  L2_31_31  5.188803e-04
K1_10_11  L1_10_10  L1_11_11  3.799708e-01
K2_10_11  L2_10_10  L2_11_11  3.799708e-01
K1_10_12  L1_10_10  L1_12_12  2.731359e-02
K2_10_12  L2_10_10  L2_12_12  2.731359e-02
K1_10_13  L1_10_10  L1_13_13  3.344225e-02
K2_10_13  L2_10_10  L2_13_13  3.344225e-02
K1_10_14  L1_10_10  L1_14_14  1.361323e-02
K2_10_14  L2_10_10  L2_14_14  1.361323e-02
K1_10_15  L1_10_10  L1_15_15  7.500458e-03
K2_10_15  L2_10_10  L2_15_15  7.500458e-03
K1_10_16  L1_10_10  L1_16_16  5.564136e-04
K2_10_16  L2_10_10  L2_16_16  5.564136e-04
K1_10_17  L1_10_10  L1_17_17  4.827563e-04
K2_10_17  L2_10_10  L2_17_17  4.827563e-04
K1_10_18  L1_10_10  L1_18_18  5.217794e-04
K2_10_18  L2_10_10  L2_18_18  5.217794e-04
K1_10_19  L1_10_10  L1_19_19  5.219556e-04
K2_10_19  L2_10_10  L2_19_19  5.219556e-04
K1_10_20  L1_10_10  L1_20_20  5.234522e-04
K2_10_20  L2_10_10  L2_20_20  5.234522e-04
K1_10_21  L1_10_10  L1_21_21  5.255776e-04
K2_10_21  L2_10_10  L2_21_21  5.255776e-04
K1_10_22  L1_10_10  L1_22_22  5.717478e-04
K2_10_22  L2_10_10  L2_22_22  5.717478e-04
K1_10_23  L1_10_10  L1_23_23  5.635897e-04
K2_10_23  L2_10_10  L2_23_23  5.635897e-04
K1_10_24  L1_10_10  L1_24_24  5.233917e-04
K2_10_24  L2_10_10  L2_24_24  5.233917e-04
K1_10_25  L1_10_10  L1_25_25  5.159250e-04
K2_10_25  L2_10_10  L2_25_25  5.159250e-04
K1_10_26  L1_10_10  L1_26_26  4.799737e-04
K2_10_26  L2_10_10  L2_26_26  4.799737e-04
K1_10_27  L1_10_10  L1_27_27  4.832980e-04
K2_10_27  L2_10_10  L2_27_27  4.832980e-04
K1_10_28  L1_10_10  L1_28_28  5.195901e-04
K2_10_28  L2_10_10  L2_28_28  5.195901e-04
K1_10_29  L1_10_10  L1_29_29  5.228041e-04
K2_10_29  L2_10_10  L2_29_29  5.228041e-04
K1_10_30  L1_10_10  L1_30_30  5.149071e-04
K2_10_30  L2_10_10  L2_30_30  5.149071e-04
K1_10_31  L1_10_10  L1_31_31  4.987550e-04
K2_10_31  L2_10_10  L2_31_31  4.987550e-04
K1_11_12  L1_11_11  L1_12_12  2.968395e-02
K2_11_12  L2_11_11  L2_12_12  2.968395e-02
K1_11_13  L1_11_11  L1_13_13  4.057717e-02
K2_11_13  L2_11_11  L2_13_13  4.057717e-02
K1_11_14  L1_11_11  L1_14_14  1.818038e-02
K2_11_14  L2_11_11  L2_14_14  1.818038e-02
K1_11_15  L1_11_11  L1_15_15  9.643380e-03
K2_11_15  L2_11_11  L2_15_15  9.643380e-03
K1_11_16  L1_11_11  L1_16_16  5.628421e-04
K2_11_16  L2_11_11  L2_16_16  5.628421e-04
K1_11_17  L1_11_11  L1_17_17  4.890381e-04
K2_11_17  L2_11_11  L2_17_17  4.890381e-04
K1_11_18  L1_11_11  L1_18_18  5.287779e-04
K2_11_18  L2_11_11  L2_18_18  5.287779e-04
K1_11_19  L1_11_11  L1_19_19  5.254044e-04
K2_11_19  L2_11_11  L2_19_19  5.254044e-04
K1_11_20  L1_11_11  L1_20_20  5.306420e-04
K2_11_20  L2_11_11  L2_20_20  5.306420e-04
K1_11_21  L1_11_11  L1_21_21  5.376005e-04
K2_11_21  L2_11_11  L2_21_21  5.376005e-04
K1_11_22  L1_11_11  L1_22_22  5.849809e-04
K2_11_22  L2_11_11  L2_22_22  5.849809e-04
K1_11_23  L1_11_11  L1_23_23  5.732865e-04
K2_11_23  L2_11_11  L2_23_23  5.732865e-04
K1_11_24  L1_11_11  L1_24_24  5.289581e-04
K2_11_24  L2_11_11  L2_24_24  5.289581e-04
K1_11_25  L1_11_11  L1_25_25  5.249464e-04
K2_11_25  L2_11_11  L2_25_25  5.249464e-04
K1_11_26  L1_11_11  L1_26_26  4.888725e-04
K2_11_26  L2_11_11  L2_26_26  4.888725e-04
K1_11_27  L1_11_11  L1_27_27  4.988859e-04
K2_11_27  L2_11_11  L2_27_27  4.988859e-04
K1_11_28  L1_11_11  L1_28_28  5.310788e-04
K2_11_28  L2_11_11  L2_28_28  5.310788e-04
K1_11_29  L1_11_11  L1_29_29  5.378607e-04
K2_11_29  L2_11_11  L2_29_29  5.378607e-04
K1_11_30  L1_11_11  L1_30_30  5.283242e-04
K2_11_30  L2_11_11  L2_30_30  5.283242e-04
K1_11_31  L1_11_11  L1_31_31  4.994429e-04
K2_11_31  L2_11_11  L2_31_31  4.994429e-04
K1_12_13  L1_12_12  L1_13_13  5.560323e-02
K2_12_13  L2_12_12  L2_13_13  5.560323e-02
K1_12_14  L1_12_12  L1_14_14  1.549013e-02
K2_12_14  L2_12_12  L2_14_14  1.549013e-02
K1_12_15  L1_12_12  L1_15_15  1.354830e-02
K2_12_15  L2_12_12  L2_15_15  1.354830e-02
K1_12_16  L1_12_12  L1_16_16  6.008719e-04
K2_12_16  L2_12_12  L2_16_16  6.008719e-04
K1_12_17  L1_12_12  L1_17_17  5.140811e-04
K2_12_17  L2_12_12  L2_17_17  5.140811e-04
K1_12_18  L1_12_12  L1_18_18  5.487191e-04
K2_12_18  L2_12_12  L2_18_18  5.487191e-04
K1_12_19  L1_12_12  L1_19_19  5.456602e-04
K2_12_19  L2_12_12  L2_19_19  5.456602e-04
K1_12_20  L1_12_12  L1_20_20  5.452295e-04
K2_12_20  L2_12_12  L2_20_20  5.452295e-04
K1_12_21  L1_12_12  L1_21_21  5.557593e-04
K2_12_21  L2_12_12  L2_21_21  5.557593e-04
K1_12_22  L1_12_12  L1_22_22  6.036344e-04
K2_12_22  L2_12_12  L2_22_22  6.036344e-04
K1_12_23  L1_12_12  L1_23_23  5.951436e-04
K2_12_23  L2_12_12  L2_23_23  5.951436e-04
K1_12_24  L1_12_12  L1_24_24  5.546356e-04
K2_12_24  L2_12_12  L2_24_24  5.546356e-04
K1_12_25  L1_12_12  L1_25_25  5.514062e-04
K2_12_25  L2_12_12  L2_25_25  5.514062e-04
K1_12_26  L1_12_12  L1_26_26  5.156899e-04
K2_12_26  L2_12_12  L2_26_26  5.156899e-04
K1_12_27  L1_12_12  L1_27_27  5.243832e-04
K2_12_27  L2_12_12  L2_27_27  5.243832e-04
K1_12_28  L1_12_12  L1_28_28  5.587464e-04
K2_12_28  L2_12_12  L2_28_28  5.587464e-04
K1_12_29  L1_12_12  L1_29_29  5.679304e-04
K2_12_29  L2_12_12  L2_29_29  5.679304e-04
K1_12_30  L1_12_12  L1_30_30  5.618144e-04
K2_12_30  L2_12_12  L2_30_30  5.618144e-04
K1_12_31  L1_12_12  L1_31_31  5.370999e-04
K2_12_31  L2_12_12  L2_31_31  5.370999e-04
K1_13_14  L1_13_13  L1_14_14  2.617642e-02
K2_13_14  L2_13_13  L2_14_14  2.617642e-02
K1_13_15  L1_13_13  L1_15_15  1.870938e-02
K2_13_15  L2_13_13  L2_15_15  1.870938e-02
K1_13_16  L1_13_13  L1_16_16  5.931027e-04
K2_13_16  L2_13_13  L2_16_16  5.931027e-04
K1_13_17  L1_13_13  L1_17_17  5.068458e-04
K2_13_17  L2_13_13  L2_17_17  5.068458e-04
K1_13_18  L1_13_13  L1_18_18  5.407514e-04
K2_13_18  L2_13_13  L2_18_18  5.407514e-04
K1_13_19  L1_13_13  L1_19_19  5.356641e-04
K2_13_19  L2_13_13  L2_19_19  5.356641e-04
K1_13_20  L1_13_13  L1_20_20  5.362053e-04
K2_13_20  L2_13_13  L2_20_20  5.362053e-04
K1_13_21  L1_13_13  L1_21_21  5.468654e-04
K2_13_21  L2_13_13  L2_21_21  5.468654e-04
K1_13_22  L1_13_13  L1_22_22  5.946096e-04
K2_13_22  L2_13_13  L2_22_22  5.946096e-04
K1_13_23  L1_13_13  L1_23_23  5.862247e-04
K2_13_23  L2_13_13  L2_23_23  5.862247e-04
K1_13_24  L1_13_13  L1_24_24  5.459538e-04
K2_13_24  L2_13_13  L2_24_24  5.459538e-04
K1_13_25  L1_13_13  L1_25_25  5.428655e-04
K2_13_25  L2_13_13  L2_25_25  5.428655e-04
K1_13_26  L1_13_13  L1_26_26  5.076389e-04
K2_13_26  L2_13_13  L2_26_26  5.076389e-04
K1_13_27  L1_13_13  L1_27_27  5.187926e-04
K2_13_27  L2_13_13  L2_27_27  5.187926e-04
K1_13_28  L1_13_13  L1_28_28  5.511800e-04
K2_13_28  L2_13_13  L2_28_28  5.511800e-04
K1_13_29  L1_13_13  L1_29_29  5.622094e-04
K2_13_29  L2_13_13  L2_29_29  5.622094e-04
K1_13_30  L1_13_13  L1_30_30  5.573657e-04
K2_13_30  L2_13_13  L2_30_30  5.573657e-04
K1_13_31  L1_13_13  L1_31_31  5.287513e-04
K2_13_31  L2_13_13  L2_31_31  5.287513e-04
K1_14_15  L1_14_14  L1_15_15  1.316875e-02
K2_14_15  L2_14_14  L2_15_15  1.316875e-02
K1_14_16  L1_14_14  L1_16_16  5.818759e-04
K2_14_16  L2_14_14  L2_16_16  5.818759e-04
K1_14_17  L1_14_14  L1_17_17  4.854675e-04
K2_14_17  L2_14_14  L2_17_17  4.854675e-04
K1_14_18  L1_14_14  L1_18_18  5.219078e-04
K2_14_18  L2_14_14  L2_18_18  5.219078e-04
K1_14_19  L1_14_14  L1_19_19  5.045642e-04
K2_14_19  L2_14_14  L2_19_19  5.045642e-04
K1_14_20  L1_14_14  L1_20_20  5.035377e-04
K2_14_20  L2_14_14  L2_20_20  5.035377e-04
K1_14_21  L1_14_14  L1_21_21  5.183612e-04
K2_14_21  L2_14_14  L2_21_21  5.183612e-04
K1_14_22  L1_14_14  L1_22_22  5.614741e-04
K2_14_22  L2_14_14  L2_22_22  5.614741e-04
K1_14_23  L1_14_14  L1_23_23  5.531796e-04
K2_14_23  L2_14_14  L2_23_23  5.531796e-04
K1_14_24  L1_14_14  L1_24_24  5.193244e-04
K2_14_24  L2_14_14  L2_24_24  5.193244e-04
K1_14_25  L1_14_14  L1_25_25  5.100664e-04
K2_14_25  L2_14_14  L2_25_25  5.100664e-04
K1_14_26  L1_14_14  L1_26_26  4.902127e-04
K2_14_26  L2_14_14  L2_26_26  4.902127e-04
K1_14_27  L1_14_14  L1_27_27  4.906665e-04
K2_14_27  L2_14_14  L2_27_27  4.906665e-04
K1_14_28  L1_14_14  L1_28_28  5.250772e-04
K2_14_28  L2_14_14  L2_28_28  5.250772e-04
K1_14_29  L1_14_14  L1_29_29  5.317526e-04
K2_14_29  L2_14_14  L2_29_29  5.317526e-04
K1_14_30  L1_14_14  L1_30_30  5.563588e-04
K2_14_30  L2_14_14  L2_30_30  5.563588e-04
K1_14_31  L1_14_14  L1_31_31  5.574840e-04
K2_14_31  L2_14_14  L2_31_31  5.574840e-04
K1_15_16  L1_15_15  L1_16_16  5.716910e-04
K2_15_16  L2_15_15  L2_16_16  5.716910e-04
K1_15_17  L1_15_15  L1_17_17  4.932378e-04
K2_15_17  L2_15_15  L2_17_17  4.932378e-04
K1_15_18  L1_15_15  L1_18_18  5.221309e-04
K2_15_18  L2_15_15  L2_18_18  5.221309e-04
K1_15_19  L1_15_15  L1_19_19  5.203094e-04
K2_15_19  L2_15_15  L2_19_19  5.203094e-04
K1_15_20  L1_15_15  L1_20_20  5.205231e-04
K2_15_20  L2_15_15  L2_20_20  5.205231e-04
K1_15_21  L1_15_15  L1_21_21  5.305933e-04
K2_15_21  L2_15_15  L2_21_21  5.305933e-04
K1_15_22  L1_15_15  L1_22_22  5.771376e-04
K2_15_22  L2_15_15  L2_22_22  5.771376e-04
K1_15_23  L1_15_15  L1_23_23  5.697039e-04
K2_15_23  L2_15_15  L2_23_23  5.697039e-04
K1_15_24  L1_15_15  L1_24_24  5.308794e-04
K2_15_24  L2_15_15  L2_24_24  5.308794e-04
K1_15_25  L1_15_15  L1_25_25  5.295346e-04
K2_15_25  L2_15_15  L2_25_25  5.295346e-04
K1_15_26  L1_15_15  L1_26_26  4.897272e-04
K2_15_26  L2_15_15  L2_26_26  4.897272e-04
K1_15_27  L1_15_15  L1_27_27  5.089421e-04
K2_15_27  L2_15_15  L2_27_27  5.089421e-04
K1_15_28  L1_15_15  L1_28_28  5.369038e-04
K2_15_28  L2_15_15  L2_28_28  5.369038e-04
K1_15_29  L1_15_15  L1_29_29  5.519604e-04
K2_15_29  L2_15_15  L2_29_29  5.519604e-04
K1_15_30  L1_15_15  L1_30_30  5.334583e-04
K2_15_30  L2_15_15  L2_30_30  5.334583e-04
K1_15_31  L1_15_15  L1_31_31  5.066535e-04
K2_15_31  L2_15_15  L2_31_31  5.066535e-04
K1_16_17  L1_16_16  L1_17_17  3.694750e-01
K2_16_17  L2_16_16  L2_17_17  3.694750e-01
K1_16_18  L1_16_16  L1_18_18  2.564489e-02
K2_16_18  L2_16_16  L2_18_18  2.564489e-02
K1_16_19  L1_16_16  L1_19_19  2.410668e-02
K2_16_19  L2_16_16  L2_19_19  2.410668e-02
K1_16_20  L1_16_16  L1_20_20  4.202120e-03
K2_16_20  L2_16_16  L2_20_20  4.202120e-03
K1_16_21  L1_16_16  L1_21_21  3.189870e-03
K2_16_21  L2_16_16  L2_21_21  3.189870e-03
K1_16_22  L1_16_16  L1_22_22  1.141627e-03
K2_16_22  L2_16_16  L2_22_22  1.141627e-03
K1_16_23  L1_16_16  L1_23_23  1.009851e-03
K2_16_23  L2_16_16  L2_23_23  1.009851e-03
K1_16_24  L1_16_16  L1_24_24  6.506150e-04
K2_16_24  L2_16_16  L2_24_24  6.506150e-04
K1_16_25  L1_16_16  L1_25_25  6.120480e-04
K2_16_25  L2_16_16  L2_25_25  6.120480e-04
K1_16_26  L1_16_16  L1_26_26  4.620545e-04
K2_16_26  L2_16_16  L2_26_26  4.620545e-04
K1_16_27  L1_16_16  L1_27_27  4.815570e-04
K2_16_27  L2_16_16  L2_27_27  4.815570e-04
K1_16_28  L1_16_16  L1_28_28  5.993057e-04
K2_16_28  L2_16_16  L2_28_28  5.993057e-04
K1_16_29  L1_16_16  L1_29_29  6.066773e-04
K2_16_29  L2_16_16  L2_29_29  6.066773e-04
K1_16_30  L1_16_16  L1_30_30  5.977872e-04
K2_16_30  L2_16_16  L2_30_30  5.977872e-04
K1_16_31  L1_16_16  L1_31_31  5.720357e-04
K2_16_31  L2_16_16  L2_31_31  5.720357e-04
K1_17_18  L1_17_17  L1_18_18  4.570846e-02
K2_17_18  L2_17_17  L2_18_18  4.570846e-02
K1_17_19  L1_17_17  L1_19_19  4.909564e-02
K2_17_19  L2_17_17  L2_19_19  4.909564e-02
K1_17_20  L1_17_17  L1_20_20  8.290244e-03
K2_17_20  L2_17_17  L2_20_20  8.290244e-03
K1_17_21  L1_17_17  L1_21_21  6.064813e-03
K2_17_21  L2_17_17  L2_21_21  6.064813e-03
K1_17_22  L1_17_17  L1_22_22  1.919467e-03
K2_17_22  L2_17_17  L2_22_22  1.919467e-03
K1_17_23  L1_17_17  L1_23_23  1.556567e-03
K2_17_23  L2_17_17  L2_23_23  1.556567e-03
K1_17_24  L1_17_17  L1_24_24  6.680015e-04
K2_17_24  L2_17_17  L2_24_24  6.680015e-04
K1_17_25  L1_17_17  L1_25_25  6.106537e-04
K2_17_25  L2_17_17  L2_25_25  6.106537e-04
K1_17_26  L1_17_17  L1_26_26  5.161500e-04
K2_17_26  L2_17_17  L2_26_26  5.161500e-04
K1_17_27  L1_17_17  L1_27_27  4.960553e-04
K2_17_27  L2_17_17  L2_27_27  4.960553e-04
K1_17_28  L1_17_17  L1_28_28  5.310886e-04
K2_17_28  L2_17_17  L2_28_28  5.310886e-04
K1_17_29  L1_17_17  L1_29_29  5.305916e-04
K2_17_29  L2_17_17  L2_29_29  5.305916e-04
K1_17_30  L1_17_17  L1_30_30  5.130697e-04
K2_17_30  L2_17_17  L2_30_30  5.130697e-04
K1_17_31  L1_17_17  L1_31_31  4.874995e-04
K2_17_31  L2_17_17  L2_31_31  4.874995e-04
K1_18_19  L1_18_18  L1_19_19  4.089782e-01
K2_18_19  L2_18_18  L2_19_19  4.089782e-01
K1_18_20  L1_18_18  L1_20_20  5.866505e-02
K2_18_20  L2_18_18  L2_20_20  5.866505e-02
K1_18_21  L1_18_18  L1_21_21  4.268254e-02
K2_18_21  L2_18_18  L2_21_21  4.268254e-02
K1_18_22  L1_18_18  L1_22_22  1.300314e-02
K2_18_22  L2_18_18  L2_22_22  1.300314e-02
K1_18_23  L1_18_18  L1_23_23  1.001745e-02
K2_18_23  L2_18_18  L2_23_23  1.001745e-02
K1_18_24  L1_18_18  L1_24_24  1.868480e-03
K2_18_24  L2_18_18  L2_24_24  1.868480e-03
K1_18_25  L1_18_18  L1_25_25  9.184351e-04
K2_18_25  L2_18_18  L2_25_25  9.184351e-04
K1_18_26  L1_18_18  L1_26_26  7.008020e-04
K2_18_26  L2_18_18  L2_26_26  7.008020e-04
K1_18_27  L1_18_18  L1_27_27  5.906962e-04
K2_18_27  L2_18_18  L2_27_27  5.906962e-04
K1_18_28  L1_18_18  L1_28_28  7.320607e-04
K2_18_28  L2_18_18  L2_28_28  7.320607e-04
K1_18_29  L1_18_18  L1_29_29  7.075982e-04
K2_18_29  L2_18_18  L2_29_29  7.075982e-04
K1_18_30  L1_18_18  L1_30_30  5.770301e-04
K2_18_30  L2_18_18  L2_30_30  5.770301e-04
K1_18_31  L1_18_18  L1_31_31  6.248162e-04
K2_18_31  L2_18_18  L2_31_31  6.248162e-04
K1_19_20  L1_19_19  L1_20_20  8.846433e-02
K2_19_20  L2_19_19  L2_20_20  8.846433e-02
K1_19_21  L1_19_19  L1_21_21  6.151794e-02
K2_19_21  L2_19_19  L2_21_21  6.151794e-02
K1_19_22  L1_19_19  L1_22_22  1.954456e-02
K2_19_22  L2_19_19  L2_22_22  1.954456e-02
K1_19_23  L1_19_19  L1_23_23  1.456527e-02
K2_19_23  L2_19_19  L2_23_23  1.456527e-02
K1_19_24  L1_19_19  L1_24_24  2.383668e-03
K2_19_24  L2_19_19  L2_24_24  2.383668e-03
K1_19_25  L1_19_19  L1_25_25  1.168580e-03
K2_19_25  L2_19_19  L2_25_25  1.168580e-03
K1_19_26  L1_19_19  L1_26_26  8.413823e-04
K2_19_26  L2_19_19  L2_26_26  8.413823e-04
K1_19_27  L1_19_19  L1_27_27  5.778551e-04
K2_19_27  L2_19_19  L2_27_27  5.778551e-04
K1_19_28  L1_19_19  L1_28_28  7.846120e-04
K2_19_28  L2_19_19  L2_28_28  7.846120e-04
K1_19_29  L1_19_19  L1_29_29  7.632200e-04
K2_19_29  L2_19_19  L2_29_29  7.632200e-04
K1_19_30  L1_19_19  L1_30_30  5.731963e-04
K2_19_30  L2_19_19  L2_30_30  5.731963e-04
K1_19_31  L1_19_19  L1_31_31  6.745317e-04
K2_19_31  L2_19_19  L2_31_31  6.745317e-04
K1_20_21  L1_20_20  L1_21_21  4.306592e-01
K2_20_21  L2_20_20  L2_21_21  4.306592e-01
K1_20_22  L1_20_20  L1_22_22  8.021498e-02
K2_20_22  L2_20_20  L2_22_22  8.021498e-02
K1_20_23  L1_20_20  L1_23_23  5.820738e-02
K2_20_23  L2_20_20  L2_23_23  5.820738e-02
K1_20_24  L1_20_20  L1_24_24  4.668546e-03
K2_20_24  L2_20_20  L2_24_24  4.668546e-03
K1_20_25  L1_20_20  L1_25_25  2.812327e-03
K2_20_25  L2_20_20  L2_25_25  2.812327e-03
K1_20_26  L1_20_20  L1_26_26  1.613459e-03
K2_20_26  L2_20_20  L2_26_26  1.613459e-03
K1_20_27  L1_20_20  L1_27_27  7.220010e-04
K2_20_27  L2_20_20  L2_27_27  7.220010e-04
K1_20_28  L1_20_20  L1_28_28  1.089887e-03
K2_20_28  L2_20_20  L2_28_28  1.089887e-03
K1_20_29  L1_20_20  L1_29_29  9.725585e-04
K2_20_29  L2_20_20  L2_29_29  9.725585e-04
K1_20_30  L1_20_20  L1_30_30  6.321237e-04
K2_20_30  L2_20_20  L2_30_30  6.321237e-04
K1_20_31  L1_20_20  L1_31_31  7.973790e-04
K2_20_31  L2_20_20  L2_31_31  7.973790e-04
K1_21_22  L1_21_21  L1_22_22  1.100919e-01
K2_21_22  L2_21_21  L2_22_22  1.100919e-01
K1_21_23  L1_21_21  L1_23_23  7.921340e-02
K2_21_23  L2_21_21  L2_23_23  7.921340e-02
K1_21_24  L1_21_21  L1_24_24  6.474059e-03
K2_21_24  L2_21_21  L2_24_24  6.474059e-03
K1_21_25  L1_21_21  L1_25_25  2.308315e-03
K2_21_25  L2_21_21  L2_25_25  2.308315e-03
K1_21_26  L1_21_21  L1_26_26  1.821661e-03
K2_21_26  L2_21_21  L2_26_26  1.821661e-03
K1_21_27  L1_21_21  L1_27_27  1.059168e-03
K2_21_27  L2_21_21  L2_27_27  1.059168e-03
K1_21_28  L1_21_21  L1_28_28  1.336246e-03
K2_21_28  L2_21_21  L2_28_28  1.336246e-03
K1_21_29  L1_21_21  L1_29_29  1.209996e-03
K2_21_29  L2_21_21  L2_29_29  1.209996e-03
K1_21_30  L1_21_21  L1_30_30  6.928026e-04
K2_21_30  L2_21_21  L2_30_30  6.928026e-04
K1_21_31  L1_21_21  L1_31_31  9.961344e-04
K2_21_31  L2_21_21  L2_31_31  9.961344e-04
K1_22_23  L1_22_22  L1_23_23  4.127477e-01
K2_22_23  L2_22_22  L2_23_23  4.127477e-01
K1_22_24  L1_22_22  L1_24_24  5.075521e-02
K2_22_24  L2_22_22  L2_24_24  5.075521e-02
K1_22_25  L1_22_22  L1_25_25  3.938330e-02
K2_22_25  L2_22_22  L2_25_25  3.938330e-02
K1_22_26  L1_22_22  L1_26_26  7.457399e-03
K2_22_26  L2_22_22  L2_26_26  7.457399e-03
K1_22_27  L1_22_22  L1_27_27  4.852878e-03
K2_22_27  L2_22_22  L2_27_27  4.852878e-03
K1_22_28  L1_22_22  L1_28_28  2.007267e-03
K2_22_28  L2_22_22  L2_28_28  2.007267e-03
K1_22_29  L1_22_22  L1_29_29  1.373906e-03
K2_22_29  L2_22_22  L2_29_29  1.373906e-03
K1_22_30  L1_22_22  L1_30_30  8.254451e-04
K2_22_30  L2_22_22  L2_30_30  8.254451e-04
K1_22_31  L1_22_22  L1_31_31  8.022536e-04
K2_22_31  L2_22_22  L2_31_31  8.022536e-04
K1_23_24  L1_23_23  L1_24_24  7.965901e-02
K2_23_24  L2_23_23  L2_24_24  7.965901e-02
K1_23_25  L1_23_23  L1_25_25  5.485515e-02
K2_23_25  L2_23_23  L2_25_25  5.485515e-02
K1_23_26  L1_23_23  L1_26_26  1.130662e-02
K2_23_26  L2_23_23  L2_26_26  1.130662e-02
K1_23_27  L1_23_23  L1_27_27  7.558274e-03
K2_23_27  L2_23_23  L2_27_27  7.558274e-03
K1_23_28  L1_23_23  L1_28_28  3.205904e-03
K2_23_28  L2_23_23  L2_28_28  3.205904e-03
K1_23_29  L1_23_23  L1_29_29  2.244951e-03
K2_23_29  L2_23_23  L2_29_29  2.244951e-03
K1_23_30  L1_23_23  L1_30_30  1.012572e-03
K2_23_30  L2_23_23  L2_30_30  1.012572e-03
K1_23_31  L1_23_23  L1_31_31  1.333191e-03
K2_23_31  L2_23_23  L2_31_31  1.333191e-03
K1_24_25  L1_24_24  L1_25_25  4.827160e-01
K2_24_25  L2_24_24  L2_25_25  4.827160e-01
K1_24_26  L1_24_24  L1_26_26  1.215932e-01
K2_24_26  L2_24_24  L2_26_26  1.215932e-01
K1_24_27  L1_24_24  L1_27_27  7.818096e-02
K2_24_27  L2_24_24  L2_27_27  7.818096e-02
K1_24_28  L1_24_24  L1_28_28  2.397309e-02
K2_24_28  L2_24_24  L2_28_28  2.397309e-02
K1_24_29  L1_24_24  L1_29_29  1.418724e-02
K2_24_29  L2_24_24  L2_29_29  1.418724e-02
K1_24_30  L1_24_24  L1_30_30  4.189989e-03
K2_24_30  L2_24_24  L2_30_30  4.189989e-03
K1_24_31  L1_24_24  L1_31_31  4.433346e-03
K2_24_31  L2_24_24  L2_31_31  4.433346e-03
K1_25_26  L1_25_25  L1_26_26  1.620293e-01
K2_25_26  L2_25_25  L2_26_26  1.620293e-01
K1_25_27  L1_25_25  L1_27_27  9.694815e-02
K2_25_27  L2_25_25  L2_27_27  9.694815e-02
K1_25_28  L1_25_25  L1_28_28  2.977385e-02
K2_25_28  L2_25_25  L2_28_28  2.977385e-02
K1_25_29  L1_25_25  L1_29_29  1.832160e-02
K2_25_29  L2_25_25  L2_29_29  1.832160e-02
K1_25_30  L1_25_25  L1_30_30  5.122981e-03
K2_25_30  L2_25_25  L2_30_30  5.122981e-03
K1_25_31  L1_25_25  L1_31_31  5.988559e-03
K2_25_31  L2_25_25  L2_31_31  5.988559e-03
K1_26_27  L1_26_26  L1_27_27  3.918531e-01
K2_26_27  L2_26_26  L2_27_27  3.918531e-01
K1_26_28  L1_26_26  L1_28_28  2.904533e-02
K2_26_28  L2_26_26  L2_28_28  2.904533e-02
K1_26_29  L1_26_26  L1_29_29  3.454705e-02
K2_26_29  L2_26_26  L2_29_29  3.454705e-02
K1_26_30  L1_26_26  L1_30_30  9.734357e-03
K2_26_30  L2_26_26  L2_30_30  9.734357e-03
K1_26_31  L1_26_26  L1_31_31  1.366183e-02
K2_26_31  L2_26_26  L2_31_31  1.366183e-02
K1_27_28  L1_27_27  L1_28_28  2.878762e-02
K2_27_28  L2_27_27  L2_28_28  2.878762e-02
K1_27_29  L1_27_27  L1_29_29  3.962567e-02
K2_27_29  L2_27_27  L2_29_29  3.962567e-02
K1_27_30  L1_27_27  L1_30_30  1.306773e-02
K2_27_30  L2_27_27  L2_30_30  1.306773e-02
K1_27_31  L1_27_27  L1_31_31  1.867102e-02
K2_27_31  L2_27_27  L2_31_31  1.867102e-02
K1_28_29  L1_28_28  L1_29_29  6.518538e-02
K2_28_29  L2_28_28  L2_29_29  6.518538e-02
K1_28_30  L1_28_28  L1_30_30  1.883694e-02
K2_28_30  L2_28_28  L2_30_30  1.883694e-02
K1_28_31  L1_28_28  L1_31_31  1.915134e-02
K2_28_31  L2_28_28  L2_31_31  1.915134e-02
K1_29_30  L1_29_29  L1_30_30  2.355387e-02
K2_29_30  L2_29_29  L2_30_30  2.355387e-02
K1_29_31  L1_29_29  L1_31_31  2.946710e-02
K2_29_31  L2_29_29  L2_31_31  2.946710e-02
K1_30_31  L1_30_30  L1_31_31  1.581045e-02
K2_30_31  L2_30_30  L2_31_31  1.581045e-02
R_G_0_0_0_0  FCHIP_RXDATA0+_Group_mid  0  1.714989e+05
C_0_0_0_0  FCHIP_RXDATA0+_Group_mid  0  3.443074e-13
R_G_1_1_1_1  FCHIP_RXDATA0-_Group_mid  0  1.667447e+05
C_1_1_1_1  FCHIP_RXDATA0-_Group_mid  0  3.542075e-13
R_G_2_2_2_2  FCHIP_RXDATA1+_Group_mid  0  1.650293e+05
C_2_2_2_2  FCHIP_RXDATA1+_Group_mid  0  3.612500e-13
R_G_3_3_3_3  FCHIP_RXDATA1-_Group_mid  0  1.776464e+05
C_3_3_3_3  FCHIP_RXDATA1-_Group_mid  0  3.258173e-13
R_G_4_4_4_4  FCHIP_RXDATA2+_Group_mid  0  1.809004e+05
C_4_4_4_4  FCHIP_RXDATA2+_Group_mid  0  3.255987e-13
R_G_5_5_5_5  FCHIP_RXDATA2-_Group_mid  0  1.886597e+05
C_5_5_5_5  FCHIP_RXDATA2-_Group_mid  0  3.030991e-13
R_G_6_6_6_6  FCHIP_RXDATA3+_Group_mid  0  2.007308e+05
C_6_6_6_6  FCHIP_RXDATA3+_Group_mid  0  2.837561e-13
R_G_7_7_7_7  FCHIP_RXDATA3-_Group_mid  0  1.954357e+05
C_7_7_7_7  FCHIP_RXDATA3-_Group_mid  0  2.936499e-13
R_G_8_8_8_8  FCHIP_RXDATA4+_Group_mid  0  1.777588e+05
C_8_8_8_8  FCHIP_RXDATA4+_Group_mid  0  3.282187e-13
R_G_9_9_9_9  FCHIP_RXDATA4-_Group_mid  0  1.810969e+05
C_9_9_9_9  FCHIP_RXDATA4-_Group_mid  0  3.207587e-13
R_G_10_10_10_10  FCHIP_RXDATA5+_Group_mid  0  1.494989e+05
C_10_10_10_10  FCHIP_RXDATA5+_Group_mid  0  4.037626e-13
R_G_11_11_11_11  FCHIP_RXDATA5-_Group_mid  0  1.494937e+05
C_11_11_11_11  FCHIP_RXDATA5-_Group_mid  0  4.033747e-13
R_G_12_12_12_12  FCHIP_RXDATA6+_Group_mid  0  1.955489e+05
C_12_12_12_12  FCHIP_RXDATA6+_Group_mid  0  2.794007e-13
R_G_13_13_13_13  FCHIP_RXDATA6-_Group_mid  0  1.929435e+05
C_13_13_13_13  FCHIP_RXDATA6-_Group_mid  0  2.829852e-13
R_G_14_14_14_14  FCHIP_RXDATA7+_Group_mid  0  1.819921e+05
C_14_14_14_14  FCHIP_RXDATA7+_Group_mid  0  3.020387e-13
R_G_15_15_15_15  FCHIP_RXDATA7-_Group_mid  0  1.876281e+05
C_15_15_15_15  FCHIP_RXDATA7-_Group_mid  0  2.922377e-13
R_G_16_16_16_16  FCHIP_TXDATA0+_Group_mid  0  1.724105e+05
C_16_16_16_16  FCHIP_TXDATA0+_Group_mid  0  3.428098e-13
R_G_17_17_17_17  FCHIP_TXDATA0-_Group_mid  0  1.661063e+05
C_17_17_17_17  FCHIP_TXDATA0-_Group_mid  0  3.575873e-13
R_G_18_18_18_18  FCHIP_TXDATA1+_Group_mid  0  1.683665e+05
C_18_18_18_18  FCHIP_TXDATA1+_Group_mid  0  3.525476e-13
R_G_19_19_19_19  FCHIP_TXDATA1-_Group_mid  0  1.651959e+05
C_19_19_19_19  FCHIP_TXDATA1-_Group_mid  0  3.608008e-13
R_G_20_20_20_20  FCHIP_TXDATA2+_Group_mid  0  1.710786e+05
C_20_20_20_20  FCHIP_TXDATA2+_Group_mid  0  3.474564e-13
R_G_21_21_21_21  FCHIP_TXDATA2-_Group_mid  0  1.760896e+05
C_21_21_21_21  FCHIP_TXDATA2-_Group_mid  0  3.322836e-13
R_G_22_22_22_22  FCHIP_TXDATA3+_Group_mid  0  1.855110e+05
C_22_22_22_22  FCHIP_TXDATA3+_Group_mid  0  3.159320e-13
R_G_23_23_23_23  FCHIP_TXDATA3-_Group_mid  0  1.950503e+05
C_23_23_23_23  FCHIP_TXDATA3-_Group_mid  0  2.939750e-13
R_G_24_24_24_24  FCHIP_TXDATA4+_Group_mid  0  1.826490e+05
C_24_24_24_24  FCHIP_TXDATA4+_Group_mid  0  3.184911e-13
R_G_25_25_25_25  FCHIP_TXDATA4-_Group_mid  0  1.816580e+05
C_25_25_25_25  FCHIP_TXDATA4-_Group_mid  0  3.203372e-13
R_G_26_26_26_26  FCHIP_TXDATA5+_Group_mid  0  1.501920e+05
C_26_26_26_26  FCHIP_TXDATA5+_Group_mid  0  4.020015e-13
R_G_27_27_27_27  FCHIP_TXDATA5-_Group_mid  0  1.493443e+05
C_27_27_27_27  FCHIP_TXDATA5-_Group_mid  0  4.038187e-13
R_G_28_28_28_28  FCHIP_TXDATA6+_Group_mid  0  1.927746e+05
C_28_28_28_28  FCHIP_TXDATA6+_Group_mid  0  2.839589e-13
R_G_29_29_29_29  FCHIP_TXDATA6-_Group_mid  0  1.924650e+05
C_29_29_29_29  FCHIP_TXDATA6-_Group_mid  0  2.836285e-13
R_G_30_30_30_30  FCHIP_TXDATA7+_Group_mid  0  1.906000e+05
C_30_30_30_30  FCHIP_TXDATA7+_Group_mid  0  2.874336e-13
R_G_31_31_31_31  FCHIP_TXDATA7-_Group_mid  0  1.830605e+05
C_31_31_31_31  FCHIP_TXDATA7-_Group_mid  0  3.002259e-13
R_G_32_32_32_32  FCHIP_VSS_Group_mid  0  1.000000e+09
C_32_32_32_32  FCHIP_VSS_Group_mid  0  1.000000e-17
C_0_1_0_1  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA0-_Group_mid  7.943466e-14
R_G_0_2_0_2  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA1+_Group_mid  8.128553e+08
C_0_2_0_2  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA1+_Group_mid  9.151865e-17
R_G_0_3_0_3  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA1-_Group_mid  1.076200e+08
C_0_3_0_3  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA1-_Group_mid  7.203267e-16
R_G_0_4_0_4  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA2+_Group_mid  1.000000e+09
C_0_4_0_4  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA2+_Group_mid  1.307248e-18
R_G_0_5_0_5  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA2-_Group_mid  1.000000e+09
C_0_5_0_5  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA2-_Group_mid  2.910317e-17
R_G_0_6_0_6  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA3+_Group_mid  1.000000e+09
C_0_6_0_6  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA3+_Group_mid  6.472047e-20
R_G_0_7_0_7  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA3-_Group_mid  1.000000e+09
C_0_7_0_7  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA3-_Group_mid  8.096630e-20
R_G_0_8_0_8  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA4+_Group_mid  1.000000e+09
C_0_8_0_8  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA4+_Group_mid  6.141825e-20
R_G_0_9_0_9  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA4-_Group_mid  1.000000e+09
C_0_9_0_9  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA4-_Group_mid  7.601717e-20
R_G_0_10_0_10  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA5+_Group_mid  1.000000e+09
C_0_10_0_10  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA5+_Group_mid  7.003276e-20
R_G_0_11_0_11  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA5-_Group_mid  1.000000e+09
C_0_11_0_11  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA5-_Group_mid  5.558149e-20
R_G_0_12_0_12  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_0_12_0_12  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA6+_Group_mid  4.965448e-20
R_G_0_13_0_13  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_0_13_0_13  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA6-_Group_mid  5.082207e-20
R_G_0_14_0_14  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_0_14_0_14  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA7+_Group_mid  5.473336e-20
R_G_0_15_0_15  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_0_15_0_15  FCHIP_RXDATA0+_Group_mid FCHIP_RXDATA7-_Group_mid  5.271276e-20
R_G_0_16_0_16  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_0_16_0_16  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA0+_Group_mid  3.243604e-20
R_G_0_17_0_17  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_0_17_0_17  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA0-_Group_mid  6.326319e-20
R_G_0_18_0_18  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_0_18_0_18  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA1+_Group_mid  5.447655e-20
R_G_0_19_0_19  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_0_19_0_19  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA1-_Group_mid  6.280633e-20
R_G_0_20_0_20  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_0_20_0_20  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA2+_Group_mid  6.077728e-20
R_G_0_21_0_21  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_0_21_0_21  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA2-_Group_mid  5.657707e-20
R_G_0_22_0_22  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_0_22_0_22  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA3+_Group_mid  5.491169e-20
R_G_0_23_0_23  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_0_23_0_23  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA3-_Group_mid  5.240107e-20
R_G_0_24_0_24  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_0_24_0_24  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA4+_Group_mid  5.541906e-20
R_G_0_25_0_25  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_0_25_0_25  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA4-_Group_mid  5.536208e-20
R_G_0_26_0_26  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_0_26_0_26  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA5+_Group_mid  7.090404e-20
R_G_0_27_0_27  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_0_27_0_27  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA5-_Group_mid  6.487966e-20
R_G_0_28_0_28  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_0_28_0_28  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA6+_Group_mid  4.728311e-20
R_G_0_29_0_29  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_0_29_0_29  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA6-_Group_mid  5.058717e-20
R_G_0_30_0_30  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_0_30_0_30  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA7+_Group_mid  5.168912e-20
R_G_0_31_0_31  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_0_31_0_31  FCHIP_RXDATA0+_Group_mid FCHIP_TXDATA7-_Group_mid  5.439221e-20
R_G_1_2_1_2  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA1+_Group_mid  1.404385e+08
C_1_2_1_2  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA1+_Group_mid  5.433943e-16
R_G_1_3_1_3  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA1-_Group_mid  4.226079e+07
C_1_3_1_3  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA1-_Group_mid  1.806042e-15
R_G_1_4_1_4  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA2+_Group_mid  1.000000e+09
C_1_4_1_4  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA2+_Group_mid  2.563657e-18
R_G_1_5_1_5  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA2-_Group_mid  1.000000e+09
C_1_5_1_5  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA2-_Group_mid  3.092341e-18
R_G_1_6_1_6  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA3+_Group_mid  1.000000e+09
C_1_6_1_6  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA3+_Group_mid  1.608714e-19
R_G_1_7_1_7  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA3-_Group_mid  1.000000e+09
C_1_7_1_7  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA3-_Group_mid  2.863602e-19
R_G_1_8_1_8  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA4+_Group_mid  1.000000e+09
C_1_8_1_8  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA4+_Group_mid  9.967124e-20
R_G_1_9_1_9  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA4-_Group_mid  1.000000e+09
C_1_9_1_9  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA4-_Group_mid  2.205754e-19
R_G_1_10_1_10  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA5+_Group_mid  1.000000e+09
C_1_10_1_10  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA5+_Group_mid  1.441102e-19
R_G_1_11_1_11  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA5-_Group_mid  1.000000e+09
C_1_11_1_11  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA5-_Group_mid  8.083452e-20
R_G_1_12_1_12  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_1_12_1_12  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA6+_Group_mid  5.171039e-20
R_G_1_13_1_13  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_1_13_1_13  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA6-_Group_mid  5.223821e-20
R_G_1_14_1_14  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_1_14_1_14  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA7+_Group_mid  5.279309e-20
R_G_1_15_1_15  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_1_15_1_15  FCHIP_RXDATA0-_Group_mid FCHIP_RXDATA7-_Group_mid  5.264525e-20
R_G_1_16_1_16  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_1_16_1_16  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA0+_Group_mid  7.081504e-20
R_G_1_17_1_17  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_1_17_1_17  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA0-_Group_mid  5.865864e-20
R_G_1_18_1_18  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_1_18_1_18  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA1+_Group_mid  5.735768e-20
R_G_1_19_1_19  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_1_19_1_19  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA1-_Group_mid  6.222354e-20
R_G_1_20_1_20  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_1_20_1_20  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA2+_Group_mid  5.119119e-20
R_G_1_21_1_21  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_1_21_1_21  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA2-_Group_mid  5.231503e-20
R_G_1_22_1_22  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_1_22_1_22  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA3+_Group_mid  5.620646e-20
R_G_1_23_1_23  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_1_23_1_23  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA3-_Group_mid  5.841278e-20
R_G_1_24_1_24  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_1_24_1_24  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA4+_Group_mid  5.181561e-20
R_G_1_25_1_25  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_1_25_1_25  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA4-_Group_mid  5.882195e-20
R_G_1_26_1_26  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_1_26_1_26  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA5+_Group_mid  7.182841e-20
R_G_1_27_1_27  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_1_27_1_27  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA5-_Group_mid  6.873279e-20
R_G_1_28_1_28  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_1_28_1_28  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA6+_Group_mid  5.589876e-20
R_G_1_29_1_29  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_1_29_1_29  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA6-_Group_mid  4.499668e-20
R_G_1_30_1_30  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_1_30_1_30  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA7+_Group_mid  4.558524e-20
R_G_1_31_1_31  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_1_31_1_31  FCHIP_RXDATA0-_Group_mid FCHIP_TXDATA7-_Group_mid  5.075735e-20
C_2_3_2_3  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA1-_Group_mid  9.043920e-14
R_G_2_4_2_4  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA2+_Group_mid  1.812691e+08
C_2_4_2_4  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA2+_Group_mid  3.904366e-16
R_G_2_5_2_5  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA2-_Group_mid  7.260603e+07
C_2_5_2_5  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA2-_Group_mid  9.334432e-16
R_G_2_6_2_6  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA3+_Group_mid  1.000000e+09
C_2_6_2_6  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA3+_Group_mid  3.362783e-19
R_G_2_7_2_7  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA3-_Group_mid  1.000000e+09
C_2_7_2_7  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA3-_Group_mid  6.447694e-19
R_G_2_8_2_8  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA4+_Group_mid  1.000000e+09
C_2_8_2_8  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA4+_Group_mid  1.646256e-19
R_G_2_9_2_9  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA4-_Group_mid  1.000000e+09
C_2_9_2_9  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA4-_Group_mid  4.577742e-19
R_G_2_10_2_10  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA5+_Group_mid  1.000000e+09
C_2_10_2_10  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA5+_Group_mid  2.529472e-19
R_G_2_11_2_11  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA5-_Group_mid  1.000000e+09
C_2_11_2_11  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA5-_Group_mid  9.454207e-20
R_G_2_12_2_12  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_2_12_2_12  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA6+_Group_mid  6.085621e-20
R_G_2_13_2_13  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_2_13_2_13  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA6-_Group_mid  6.323639e-20
R_G_2_14_2_14  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_2_14_2_14  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA7+_Group_mid  6.056859e-20
R_G_2_15_2_15  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_2_15_2_15  FCHIP_RXDATA1+_Group_mid FCHIP_RXDATA7-_Group_mid  5.784062e-20
R_G_2_16_2_16  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_2_16_2_16  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA0+_Group_mid  5.991298e-20
R_G_2_17_2_17  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_2_17_2_17  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA0-_Group_mid  5.774947e-20
R_G_2_18_2_18  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_2_18_2_18  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA1+_Group_mid  7.068082e-20
R_G_2_19_2_19  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_2_19_2_19  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA1-_Group_mid  6.601055e-20
R_G_2_20_2_20  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_2_20_2_20  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA2+_Group_mid  6.565134e-20
R_G_2_21_2_21  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_2_21_2_21  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA2-_Group_mid  6.286094e-20
R_G_2_22_2_22  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_2_22_2_22  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA3+_Group_mid  6.020299e-20
R_G_2_23_2_23  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_2_23_2_23  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA3-_Group_mid  5.857163e-20
R_G_2_24_2_24  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_2_24_2_24  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA4+_Group_mid  6.504434e-20
R_G_2_25_2_25  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_2_25_2_25  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA4-_Group_mid  6.183977e-20
R_G_2_26_2_26  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_2_26_2_26  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA5+_Group_mid  7.700384e-20
R_G_2_27_2_27  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_2_27_2_27  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA5-_Group_mid  7.329991e-20
R_G_2_28_2_28  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_2_28_2_28  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA6+_Group_mid  5.607202e-20
R_G_2_29_2_29  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_2_29_2_29  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA6-_Group_mid  5.100490e-20
R_G_2_30_2_30  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_2_30_2_30  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA7+_Group_mid  5.528295e-20
R_G_2_31_2_31  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_2_31_2_31  FCHIP_RXDATA1+_Group_mid FCHIP_TXDATA7-_Group_mid  5.532874e-20
R_G_3_4_3_4  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA2+_Group_mid  3.759485e+08
C_3_4_3_4  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA2+_Group_mid  2.191416e-16
R_G_3_5_3_5  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA2-_Group_mid  1.051437e+08
C_3_5_3_5  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA2-_Group_mid  7.435891e-16
R_G_3_6_3_6  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA3+_Group_mid  1.000000e+09
C_3_6_3_6  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA3+_Group_mid  1.900245e-19
R_G_3_7_3_7  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA3-_Group_mid  1.000000e+09
C_3_7_3_7  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA3-_Group_mid  3.497844e-19
R_G_3_8_3_8  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA4+_Group_mid  1.000000e+09
C_3_8_3_8  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA4+_Group_mid  1.073980e-19
R_G_3_9_3_9  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA4-_Group_mid  1.000000e+09
C_3_9_3_9  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA4-_Group_mid  2.564376e-19
R_G_3_10_3_10  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA5+_Group_mid  1.000000e+09
C_3_10_3_10  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA5+_Group_mid  1.604355e-19
R_G_3_11_3_11  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA5-_Group_mid  1.000000e+09
C_3_11_3_11  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA5-_Group_mid  7.643936e-20
R_G_3_12_3_12  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_3_12_3_12  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA6+_Group_mid  5.156052e-20
R_G_3_13_3_13  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_3_13_3_13  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA6-_Group_mid  5.286533e-20
R_G_3_14_3_14  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_3_14_3_14  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA7+_Group_mid  5.489278e-20
R_G_3_15_3_15  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_3_15_3_15  FCHIP_RXDATA1-_Group_mid FCHIP_RXDATA7-_Group_mid  5.015831e-20
R_G_3_16_3_16  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_3_16_3_16  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA0+_Group_mid  5.692469e-20
R_G_3_17_3_17  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_3_17_3_17  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA0-_Group_mid  4.877495e-20
R_G_3_18_3_18  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_3_18_3_18  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA1+_Group_mid  5.401869e-20
R_G_3_19_3_19  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_3_19_3_19  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA1-_Group_mid  5.741309e-20
R_G_3_20_3_20  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_3_20_3_20  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA2+_Group_mid  5.371027e-20
R_G_3_21_3_21  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_3_21_3_21  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA2-_Group_mid  5.648776e-20
R_G_3_22_3_22  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_3_22_3_22  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA3+_Group_mid  5.508945e-20
R_G_3_23_3_23  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_3_23_3_23  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA3-_Group_mid  4.810098e-20
R_G_3_24_3_24  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_3_24_3_24  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA4+_Group_mid  5.262871e-20
R_G_3_25_3_25  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_3_25_3_25  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA4-_Group_mid  5.479017e-20
R_G_3_26_3_26  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_3_26_3_26  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA5+_Group_mid  6.785950e-20
R_G_3_27_3_27  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_3_27_3_27  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA5-_Group_mid  6.337624e-20
R_G_3_28_3_28  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_3_28_3_28  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA6+_Group_mid  5.342128e-20
R_G_3_29_3_29  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_3_29_3_29  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA6-_Group_mid  4.706248e-20
R_G_3_30_3_30  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_3_30_3_30  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA7+_Group_mid  4.910010e-20
R_G_3_31_3_31  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_3_31_3_31  FCHIP_RXDATA1-_Group_mid FCHIP_TXDATA7-_Group_mid  5.049429e-20
C_4_5_4_5  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA2-_Group_mid  8.227007e-14
R_G_4_6_4_6  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA3+_Group_mid  1.846636e+08
C_4_6_4_6  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA3+_Group_mid  4.278906e-16
R_G_4_7_4_7  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA3-_Group_mid  1.003894e+08
C_4_7_4_7  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA3-_Group_mid  7.010999e-16
R_G_4_8_4_8  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA4+_Group_mid  1.000000e+09
C_4_8_4_8  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA4+_Group_mid  4.230211e-17
R_G_4_9_4_9  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA4-_Group_mid  1.000000e+09
C_4_9_4_9  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA4-_Group_mid  1.039900e-16
R_G_4_10_4_10  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA5+_Group_mid  1.000000e+09
C_4_10_4_10  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA5+_Group_mid  6.366065e-18
R_G_4_11_4_11  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA5-_Group_mid  1.000000e+09
C_4_11_4_11  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA5-_Group_mid  5.252500e-18
R_G_4_12_4_12  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_4_12_4_12  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA6+_Group_mid  6.056370e-20
R_G_4_13_4_13  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_4_13_4_13  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA6-_Group_mid  6.311896e-20
R_G_4_14_4_14  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_4_14_4_14  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA7+_Group_mid  5.950157e-20
R_G_4_15_4_15  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_4_15_4_15  FCHIP_RXDATA2+_Group_mid FCHIP_RXDATA7-_Group_mid  5.324959e-20
R_G_4_16_4_16  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_4_16_4_16  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA0+_Group_mid  5.850847e-20
R_G_4_17_4_17  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_4_17_4_17  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA0-_Group_mid  4.940347e-20
R_G_4_18_4_18  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_4_18_4_18  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA1+_Group_mid  5.841356e-20
R_G_4_19_4_19  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_4_19_4_19  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA1-_Group_mid  5.872879e-20
R_G_4_20_4_20  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_4_20_4_20  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA2+_Group_mid  5.638025e-20
R_G_4_21_4_21  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_4_21_4_21  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA2-_Group_mid  5.160841e-20
R_G_4_22_4_22  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_4_22_4_22  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA3+_Group_mid  5.298750e-20
R_G_4_23_4_23  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_4_23_4_23  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA3-_Group_mid  4.847506e-20
R_G_4_24_4_24  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_4_24_4_24  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA4+_Group_mid  5.207825e-20
R_G_4_25_4_25  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_4_25_4_25  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA4-_Group_mid  5.450390e-20
R_G_4_26_4_26  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_4_26_4_26  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA5+_Group_mid  6.793425e-20
R_G_4_27_4_27  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_4_27_4_27  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA5-_Group_mid  6.434537e-20
R_G_4_28_4_28  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_4_28_4_28  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA6+_Group_mid  4.850779e-20
R_G_4_29_4_29  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_4_29_4_29  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA6-_Group_mid  4.331166e-20
R_G_4_30_4_30  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_4_30_4_30  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA7+_Group_mid  4.879636e-20
R_G_4_31_4_31  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_4_31_4_31  FCHIP_RXDATA2+_Group_mid FCHIP_TXDATA7-_Group_mid  4.947574e-20
R_G_5_6_5_6  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA3+_Group_mid  3.471147e+08
C_5_6_5_6  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA3+_Group_mid  2.783329e-16
R_G_5_7_5_7  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA3-_Group_mid  1.800965e+08
C_5_7_5_7  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA3-_Group_mid  4.529756e-16
R_G_5_8_5_8  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA4+_Group_mid  1.000000e+09
C_5_8_5_8  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA4+_Group_mid  3.774820e-17
R_G_5_9_5_9  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA4-_Group_mid  1.000000e+09
C_5_9_5_9  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA4-_Group_mid  7.632165e-17
R_G_5_10_5_10  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA5+_Group_mid  1.000000e+09
C_5_10_5_10  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA5+_Group_mid  7.066050e-18
R_G_5_11_5_11  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA5-_Group_mid  1.000000e+09
C_5_11_5_11  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA5-_Group_mid  5.882899e-18
R_G_5_12_5_12  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_5_12_5_12  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA6+_Group_mid  5.088040e-20
R_G_5_13_5_13  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_5_13_5_13  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA6-_Group_mid  5.209311e-20
R_G_5_14_5_14  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_5_14_5_14  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA7+_Group_mid  5.246553e-20
R_G_5_15_5_15  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_5_15_5_15  FCHIP_RXDATA2-_Group_mid FCHIP_RXDATA7-_Group_mid  4.817658e-20
R_G_5_16_5_16  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_5_16_5_16  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA0+_Group_mid  5.259710e-20
R_G_5_17_5_17  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_5_17_5_17  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA0-_Group_mid  4.578996e-20
R_G_5_18_5_18  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_5_18_5_18  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA1+_Group_mid  5.535066e-20
R_G_5_19_5_19  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_5_19_5_19  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA1-_Group_mid  5.420165e-20
R_G_5_20_5_20  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_5_20_5_20  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA2+_Group_mid  5.475426e-20
R_G_5_21_5_21  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_5_21_5_21  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA2-_Group_mid  5.396016e-20
R_G_5_22_5_22  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_5_22_5_22  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA3+_Group_mid  5.346126e-20
R_G_5_23_5_23  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_5_23_5_23  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA3-_Group_mid  4.442435e-20
R_G_5_24_5_24  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_5_24_5_24  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA4+_Group_mid  5.054044e-20
R_G_5_25_5_25  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_5_25_5_25  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA4-_Group_mid  5.278995e-20
R_G_5_26_5_26  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_5_26_5_26  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA5+_Group_mid  6.435966e-20
R_G_5_27_5_27  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_5_27_5_27  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA5-_Group_mid  6.085696e-20
R_G_5_28_5_28  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_5_28_5_28  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA6+_Group_mid  5.052695e-20
R_G_5_29_5_29  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_5_29_5_29  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA6-_Group_mid  4.366494e-20
R_G_5_30_5_30  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_5_30_5_30  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA7+_Group_mid  4.717311e-20
R_G_5_31_5_31  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_5_31_5_31  FCHIP_RXDATA2-_Group_mid FCHIP_TXDATA7-_Group_mid  4.719535e-20
R_G_6_7_6_7  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA3-_Group_mid  1.048570e+06
C_6_7_6_7  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA3-_Group_mid  7.323332e-14
R_G_6_8_6_8  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA4+_Group_mid  2.580500e+07
C_6_8_6_8  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA4+_Group_mid  2.627505e-15
R_G_6_9_6_9  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA4-_Group_mid  6.900657e+06
C_6_9_6_9  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA4-_Group_mid  1.046240e-14
R_G_6_10_6_10  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA5+_Group_mid  1.000000e+09
C_6_10_6_10  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA5+_Group_mid  1.034386e-16
R_G_6_11_6_11  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA5-_Group_mid  1.000000e+09
C_6_11_6_11  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA5-_Group_mid  6.660427e-17
R_G_6_12_6_12  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_6_12_6_12  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA6+_Group_mid  5.622706e-20
R_G_6_13_6_13  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_6_13_6_13  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA6-_Group_mid  7.797924e-20
R_G_6_14_6_14  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_6_14_6_14  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA7+_Group_mid  7.202060e-20
R_G_6_15_6_15  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_6_15_6_15  FCHIP_RXDATA3+_Group_mid FCHIP_RXDATA7-_Group_mid  4.909710e-20
R_G_6_16_6_16  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_6_16_6_16  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA0+_Group_mid  4.846036e-20
R_G_6_17_6_17  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_6_17_6_17  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA0-_Group_mid  4.916621e-20
R_G_6_18_6_18  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_6_18_6_18  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA1+_Group_mid  5.046441e-20
R_G_6_19_6_19  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_6_19_6_19  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA1-_Group_mid  5.094044e-20
R_G_6_20_6_20  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_6_20_6_20  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA2+_Group_mid  5.363142e-20
R_G_6_21_6_21  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_6_21_6_21  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA2-_Group_mid  4.831520e-20
R_G_6_22_6_22  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_6_22_6_22  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA3+_Group_mid  4.554212e-20
R_G_6_23_6_23  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_6_23_6_23  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA3-_Group_mid  4.247536e-20
R_G_6_24_6_24  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_6_24_6_24  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA4+_Group_mid  5.000750e-20
R_G_6_25_6_25  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_6_25_6_25  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA4-_Group_mid  4.669240e-20
R_G_6_26_6_26  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_6_26_6_26  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA5+_Group_mid  5.996732e-20
R_G_6_27_6_27  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_6_27_6_27  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA5-_Group_mid  5.575545e-20
R_G_6_28_6_28  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_6_28_6_28  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA6+_Group_mid  4.648586e-20
R_G_6_29_6_29  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_6_29_6_29  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA6-_Group_mid  3.998240e-20
R_G_6_30_6_30  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_6_30_6_30  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA7+_Group_mid  4.394136e-20
R_G_6_31_6_31  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_6_31_6_31  FCHIP_RXDATA3+_Group_mid FCHIP_TXDATA7-_Group_mid  4.398896e-20
R_G_7_8_7_8  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA4+_Group_mid  6.564903e+07
C_7_8_7_8  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA4+_Group_mid  1.111911e-15
R_G_7_9_7_9  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA4-_Group_mid  2.391535e+07
C_7_9_7_9  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA4-_Group_mid  2.854149e-15
R_G_7_10_7_10  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA5+_Group_mid  1.000000e+09
C_7_10_7_10  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA5+_Group_mid  6.537155e-17
R_G_7_11_7_11  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA5-_Group_mid  1.000000e+09
C_7_11_7_11  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA5-_Group_mid  4.568659e-17
R_G_7_12_7_12  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_7_12_7_12  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA6+_Group_mid  4.633812e-20
R_G_7_13_7_13  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_7_13_7_13  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA6-_Group_mid  5.021592e-20
R_G_7_14_7_14  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_7_14_7_14  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA7+_Group_mid  5.132156e-20
R_G_7_15_7_15  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_7_15_7_15  FCHIP_RXDATA3-_Group_mid FCHIP_RXDATA7-_Group_mid  4.669837e-20
R_G_7_16_7_16  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_7_16_7_16  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA0+_Group_mid  5.142046e-20
R_G_7_17_7_17  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_7_17_7_17  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA0-_Group_mid  4.666522e-20
R_G_7_18_7_18  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_7_18_7_18  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA1+_Group_mid  5.255622e-20
R_G_7_19_7_19  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_7_19_7_19  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA1-_Group_mid  5.300285e-20
R_G_7_20_7_20  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_7_20_7_20  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA2+_Group_mid  5.117012e-20
R_G_7_21_7_21  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_7_21_7_21  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA2-_Group_mid  4.924094e-20
R_G_7_22_7_22  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_7_22_7_22  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA3+_Group_mid  5.000831e-20
R_G_7_23_7_23  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_7_23_7_23  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA3-_Group_mid  4.294724e-20
R_G_7_24_7_24  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_7_24_7_24  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA4+_Group_mid  4.811754e-20
R_G_7_25_7_25  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_7_25_7_25  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA4-_Group_mid  4.913321e-20
R_G_7_26_7_26  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_7_26_7_26  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA5+_Group_mid  6.150852e-20
R_G_7_27_7_27  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_7_27_7_27  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA5-_Group_mid  5.778811e-20
R_G_7_28_7_28  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_7_28_7_28  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA6+_Group_mid  3.920398e-20
R_G_7_29_7_29  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_7_29_7_29  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA6-_Group_mid  4.395879e-20
R_G_7_30_7_30  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_7_30_7_30  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA7+_Group_mid  4.425933e-20
R_G_7_31_7_31  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_7_31_7_31  FCHIP_RXDATA3-_Group_mid FCHIP_TXDATA7-_Group_mid  4.511532e-20
C_8_9_8_9  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA4-_Group_mid  8.932430e-14
R_G_8_10_8_10  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA5+_Group_mid  4.895484e+07
C_8_10_8_10  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA5+_Group_mid  1.429374e-15
R_G_8_11_8_11  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA5-_Group_mid  1.016464e+08
C_8_11_8_11  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA5-_Group_mid  7.538901e-16
R_G_8_12_8_12  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_8_12_8_12  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA6+_Group_mid  3.801485e-19
R_G_8_13_8_13  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_8_13_8_13  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA6-_Group_mid  2.918294e-19
R_G_8_14_8_14  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_8_14_8_14  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA7+_Group_mid  1.786540e-19
R_G_8_15_8_15  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_8_15_8_15  FCHIP_RXDATA4+_Group_mid FCHIP_RXDATA7-_Group_mid  1.058873e-19
R_G_8_16_8_16  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_8_16_8_16  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA0+_Group_mid  5.823495e-20
R_G_8_17_8_17  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_8_17_8_17  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA0-_Group_mid  5.453070e-20
R_G_8_18_8_18  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_8_18_8_18  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA1+_Group_mid  5.877365e-20
R_G_8_19_8_19  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_8_19_8_19  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA1-_Group_mid  5.919577e-20
R_G_8_20_8_20  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_8_20_8_20  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA2+_Group_mid  5.786458e-20
R_G_8_21_8_21  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_8_21_8_21  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA2-_Group_mid  5.539337e-20
R_G_8_22_8_22  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_8_22_8_22  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA3+_Group_mid  5.391538e-20
R_G_8_23_8_23  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_8_23_8_23  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA3-_Group_mid  5.009612e-20
R_G_8_24_8_24  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_8_24_8_24  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA4+_Group_mid  5.511830e-20
R_G_8_25_8_25  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_8_25_8_25  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA4-_Group_mid  5.456898e-20
R_G_8_26_8_26  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_8_26_8_26  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA5+_Group_mid  6.924675e-20
R_G_8_27_8_27  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_8_27_8_27  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA5-_Group_mid  6.455371e-20
R_G_8_28_8_28  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_8_28_8_28  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA6+_Group_mid  4.911160e-20
R_G_8_29_8_29  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_8_29_8_29  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA6-_Group_mid  4.849578e-20
R_G_8_30_8_30  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_8_30_8_30  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA7+_Group_mid  4.999141e-20
R_G_8_31_8_31  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_8_31_8_31  FCHIP_RXDATA4+_Group_mid FCHIP_TXDATA7-_Group_mid  5.090457e-20
R_G_9_10_9_10  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA5+_Group_mid  1.145988e+08
C_9_10_9_10  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA5+_Group_mid  6.610271e-16
R_G_9_11_9_11  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA5-_Group_mid  2.287792e+08
C_9_11_9_11  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA5-_Group_mid  3.768922e-16
R_G_9_12_9_12  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_9_12_9_12  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA6+_Group_mid  2.449223e-19
R_G_9_13_9_13  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_9_13_9_13  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA6-_Group_mid  1.966186e-19
R_G_9_14_9_14  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_9_14_9_14  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA7+_Group_mid  1.229442e-19
R_G_9_15_9_15  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_9_15_9_15  FCHIP_RXDATA4-_Group_mid FCHIP_RXDATA7-_Group_mid  8.128949e-20
R_G_9_16_9_16  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_9_16_9_16  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA0+_Group_mid  5.633848e-20
R_G_9_17_9_17  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_9_17_9_17  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA0-_Group_mid  5.283698e-20
R_G_9_18_9_18  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_9_18_9_18  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA1+_Group_mid  5.568091e-20
R_G_9_19_9_19  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_9_19_9_19  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA1-_Group_mid  5.774540e-20
R_G_9_20_9_20  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_9_20_9_20  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA2+_Group_mid  5.497973e-20
R_G_9_21_9_21  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_9_21_9_21  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA2-_Group_mid  5.748830e-20
R_G_9_22_9_22  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_9_22_9_22  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA3+_Group_mid  5.241750e-20
R_G_9_23_9_23  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_9_23_9_23  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA3-_Group_mid  4.927722e-20
R_G_9_24_9_24  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_9_24_9_24  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA4+_Group_mid  5.408118e-20
R_G_9_25_9_25  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_9_25_9_25  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA4-_Group_mid  5.307387e-20
R_G_9_26_9_26  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_9_26_9_26  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA5+_Group_mid  6.850703e-20
R_G_9_27_9_27  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_9_27_9_27  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA5-_Group_mid  6.255318e-20
R_G_9_28_9_28  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_9_28_9_28  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA6+_Group_mid  4.604790e-20
R_G_9_29_9_29  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_9_29_9_29  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA6-_Group_mid  4.846060e-20
R_G_9_30_9_30  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_9_30_9_30  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA7+_Group_mid  4.931378e-20
R_G_9_31_9_31  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_9_31_9_31  FCHIP_RXDATA4-_Group_mid FCHIP_TXDATA7-_Group_mid  4.983617e-20
C_10_11_10_11  FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA5-_Group_mid  1.156590e-13
R_G_10_12_10_12  FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_10_12_10_12  FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA6+_Group_mid  4.086136e-19
R_G_10_13_10_13  FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_10_13_10_13  FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA6-_Group_mid  7.907616e-19
R_G_10_14_10_14  FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_10_14_10_14  FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA7+_Group_mid  4.431046e-19
R_G_10_15_10_15  FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_10_15_10_15  FCHIP_RXDATA5+_Group_mid FCHIP_RXDATA7-_Group_mid  2.121858e-19
R_G_10_16_10_16  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_10_16_10_16  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA0+_Group_mid  7.342099e-20
R_G_10_17_10_17  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_10_17_10_17  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA0-_Group_mid  6.699003e-20
R_G_10_18_10_18  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_10_18_10_18  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA1+_Group_mid  7.212129e-20
R_G_10_19_10_19  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_10_19_10_19  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA1-_Group_mid  7.556691e-20
R_G_10_20_10_20  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_10_20_10_20  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA2+_Group_mid  7.340394e-20
R_G_10_21_10_21  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_10_21_10_21  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA2-_Group_mid  6.959054e-20
R_G_10_22_10_22  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_10_22_10_22  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA3+_Group_mid  6.651674e-20
R_G_10_23_10_23  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_10_23_10_23  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA3-_Group_mid  6.194633e-20
R_G_10_24_10_24  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_10_24_10_24  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA4+_Group_mid  6.739920e-20
R_G_10_25_10_25  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_10_25_10_25  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA4-_Group_mid  6.768826e-20
R_G_10_26_10_26  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_10_26_10_26  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA5+_Group_mid  8.624036e-20
R_G_10_27_10_27  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_10_27_10_27  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA5-_Group_mid  7.931582e-20
R_G_10_28_10_28  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_10_28_10_28  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA6+_Group_mid  5.998613e-20
R_G_10_29_10_29  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_10_29_10_29  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA6-_Group_mid  5.979121e-20
R_G_10_30_10_30  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_10_30_10_30  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA7+_Group_mid  6.116158e-20
R_G_10_31_10_31  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_10_31_10_31  FCHIP_RXDATA5+_Group_mid FCHIP_TXDATA7-_Group_mid  6.467108e-20
R_G_11_12_11_12  FCHIP_RXDATA5-_Group_mid FCHIP_RXDATA6+_Group_mid  1.000000e+09
C_11_12_11_12  FCHIP_RXDATA5-_Group_mid FCHIP_RXDATA6+_Group_mid  7.826934e-19
R_G_11_13_11_13  FCHIP_RXDATA5-_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_11_13_11_13  FCHIP_RXDATA5-_Group_mid FCHIP_RXDATA6-_Group_mid  1.229025e-18
R_G_11_14_11_14  FCHIP_RXDATA5-_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_11_14_11_14  FCHIP_RXDATA5-_Group_mid FCHIP_RXDATA7+_Group_mid  7.399413e-19
R_G_11_15_11_15  FCHIP_RXDATA5-_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_11_15_11_15  FCHIP_RXDATA5-_Group_mid FCHIP_RXDATA7-_Group_mid  3.742128e-19
R_G_11_16_11_16  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_11_16_11_16  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA0+_Group_mid  6.734678e-20
R_G_11_17_11_17  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_11_17_11_17  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA0-_Group_mid  6.141715e-20
R_G_11_18_11_18  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_11_18_11_18  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA1+_Group_mid  6.662404e-20
R_G_11_19_11_19  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_11_19_11_19  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA1-_Group_mid  6.950186e-20
R_G_11_20_11_20  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_11_20_11_20  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA2+_Group_mid  6.782673e-20
R_G_11_21_11_21  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_11_21_11_21  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA2-_Group_mid  6.555883e-20
R_G_11_22_11_22  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_11_22_11_22  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA3+_Group_mid  6.275167e-20
R_G_11_23_11_23  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_11_23_11_23  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA3-_Group_mid  5.783676e-20
R_G_11_24_11_24  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_11_24_11_24  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA4+_Group_mid  6.185564e-20
R_G_11_25_11_25  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_11_25_11_25  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA4-_Group_mid  6.393854e-20
R_G_11_26_11_26  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_11_26_11_26  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA5+_Group_mid  7.991833e-20
R_G_11_27_11_27  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_11_27_11_27  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA5-_Group_mid  7.564847e-20
R_G_11_28_11_28  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_11_28_11_28  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA6+_Group_mid  5.613251e-20
R_G_11_29_11_29  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_11_29_11_29  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA6-_Group_mid  5.607051e-20
R_G_11_30_11_30  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_11_30_11_30  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA7+_Group_mid  5.699686e-20
R_G_11_31_11_31  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_11_31_11_31  FCHIP_RXDATA5-_Group_mid FCHIP_TXDATA7-_Group_mid  5.771321e-20
R_G_12_13_12_13  FCHIP_RXDATA6+_Group_mid FCHIP_RXDATA6-_Group_mid  1.000000e+09
C_12_13_12_13  FCHIP_RXDATA6+_Group_mid FCHIP_RXDATA6-_Group_mid  1.044890e-18
R_G_12_14_12_14  FCHIP_RXDATA6+_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_12_14_12_14  FCHIP_RXDATA6+_Group_mid FCHIP_RXDATA7+_Group_mid  3.605707e-19
R_G_12_15_12_15  FCHIP_RXDATA6+_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_12_15_12_15  FCHIP_RXDATA6+_Group_mid FCHIP_RXDATA7-_Group_mid  2.930166e-19
R_G_12_16_12_16  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_12_16_12_16  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA0+_Group_mid  4.957354e-20
R_G_12_17_12_17  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_12_17_12_17  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA0-_Group_mid  4.543439e-20
R_G_12_18_12_18  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_12_18_12_18  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA1+_Group_mid  4.899314e-20
R_G_12_19_12_19  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_12_19_12_19  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA1-_Group_mid  5.002444e-20
R_G_12_20_12_20  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_12_20_12_20  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA2+_Group_mid  4.892578e-20
R_G_12_21_12_21  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_12_21_12_21  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA2-_Group_mid  4.776746e-20
R_G_12_22_12_22  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_12_22_12_22  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA3+_Group_mid  4.540246e-20
R_G_12_23_12_23  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_12_23_12_23  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA3-_Group_mid  4.204431e-20
R_G_12_24_12_24  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_12_24_12_24  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA4+_Group_mid  4.571232e-20
R_G_12_25_12_25  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_12_25_12_25  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA4-_Group_mid  4.609281e-20
R_G_12_26_12_26  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_12_26_12_26  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA5+_Group_mid  5.855391e-20
R_G_12_27_12_27  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_12_27_12_27  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA5-_Group_mid  5.460321e-20
R_G_12_28_12_28  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_12_28_12_28  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA6+_Group_mid  4.063406e-20
R_G_12_29_12_29  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_12_29_12_29  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA6-_Group_mid  4.087531e-20
R_G_12_30_12_30  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_12_30_12_30  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA7+_Group_mid  4.153076e-20
R_G_12_31_12_31  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_12_31_12_31  FCHIP_RXDATA6+_Group_mid FCHIP_TXDATA7-_Group_mid  4.316360e-20
R_G_13_14_13_14  FCHIP_RXDATA6-_Group_mid FCHIP_RXDATA7+_Group_mid  1.000000e+09
C_13_14_13_14  FCHIP_RXDATA6-_Group_mid FCHIP_RXDATA7+_Group_mid  6.073473e-19
R_G_13_15_13_15  FCHIP_RXDATA6-_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_13_15_13_15  FCHIP_RXDATA6-_Group_mid FCHIP_RXDATA7-_Group_mid  4.088104e-19
R_G_13_16_13_16  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_13_16_13_16  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA0+_Group_mid  5.030545e-20
R_G_13_17_13_17  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_13_17_13_17  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA0-_Group_mid  4.610643e-20
R_G_13_18_13_18  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_13_18_13_18  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA1+_Group_mid  4.983324e-20
R_G_13_19_13_19  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_13_19_13_19  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA1-_Group_mid  5.066769e-20
R_G_13_20_13_20  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_13_20_13_20  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA2+_Group_mid  4.968160e-20
R_G_13_21_13_21  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_13_21_13_21  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA2-_Group_mid  4.864513e-20
R_G_13_22_13_22  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_13_22_13_22  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA3+_Group_mid  4.612796e-20
R_G_13_23_13_23  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_13_23_13_23  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA3-_Group_mid  4.287720e-20
R_G_13_24_13_24  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_13_24_13_24  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA4+_Group_mid  4.639396e-20
R_G_13_25_13_25  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_13_25_13_25  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA4-_Group_mid  4.678069e-20
R_G_13_26_13_26  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_13_26_13_26  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA5+_Group_mid  5.932115e-20
R_G_13_27_13_27  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_13_27_13_27  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA5-_Group_mid  5.560744e-20
R_G_13_28_13_28  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_13_28_13_28  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA6+_Group_mid  4.135921e-20
R_G_13_29_13_29  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_13_29_13_29  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA6-_Group_mid  4.152555e-20
R_G_13_30_13_30  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_13_30_13_30  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA7+_Group_mid  4.228639e-20
R_G_13_31_13_31  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_13_31_13_31  FCHIP_RXDATA6-_Group_mid FCHIP_TXDATA7-_Group_mid  4.359656e-20
R_G_14_15_14_15  FCHIP_RXDATA7+_Group_mid FCHIP_RXDATA7-_Group_mid  1.000000e+09
C_14_15_14_15  FCHIP_RXDATA7+_Group_mid FCHIP_RXDATA7-_Group_mid  3.346198e-19
R_G_14_16_14_16  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_14_16_14_16  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA0+_Group_mid  5.576349e-20
R_G_14_17_14_17  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_14_17_14_17  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA0-_Group_mid  4.943325e-20
R_G_14_18_14_18  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_14_18_14_18  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA1+_Group_mid  5.680490e-20
R_G_14_19_14_19  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_14_19_14_19  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA1-_Group_mid  5.408854e-20
R_G_14_20_14_20  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_14_20_14_20  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA2+_Group_mid  5.273658e-20
R_G_14_21_14_21  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_14_21_14_21  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA2-_Group_mid  5.285525e-20
R_G_14_22_14_22  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_14_22_14_22  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA3+_Group_mid  4.940628e-20
R_G_14_23_14_23  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_14_23_14_23  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA3-_Group_mid  4.580915e-20
R_G_14_24_14_24  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_14_24_14_24  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA4+_Group_mid  5.027193e-20
R_G_14_25_14_25  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_14_25_14_25  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA4-_Group_mid  4.957795e-20
R_G_14_26_14_26  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_14_26_14_26  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA5+_Group_mid  6.502683e-20
R_G_14_27_14_27  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_14_27_14_27  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA5-_Group_mid  5.874914e-20
R_G_14_28_14_28  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_14_28_14_28  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA6+_Group_mid  4.746551e-20
R_G_14_29_14_29  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_14_29_14_29  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA6-_Group_mid  4.220144e-20
R_G_14_30_14_30  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_14_30_14_30  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA7+_Group_mid  4.681600e-20
R_G_14_31_14_31  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_14_31_14_31  FCHIP_RXDATA7+_Group_mid FCHIP_TXDATA7-_Group_mid  5.140747e-20
R_G_15_16_15_16  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA0+_Group_mid  1.000000e+09
C_15_16_15_16  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA0+_Group_mid  5.134642e-20
R_G_15_17_15_17  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA0-_Group_mid  1.000000e+09
C_15_17_15_17  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA0-_Group_mid  4.791375e-20
R_G_15_18_15_18  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA1+_Group_mid  1.000000e+09
C_15_18_15_18  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA1+_Group_mid  5.041453e-20
R_G_15_19_15_19  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_15_19_15_19  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA1-_Group_mid  5.270494e-20
R_G_15_20_15_20  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_15_20_15_20  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA2+_Group_mid  5.190691e-20
R_G_15_21_15_21  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_15_21_15_21  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA2-_Group_mid  4.950555e-20
R_G_15_22_15_22  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_15_22_15_22  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA3+_Group_mid  4.811714e-20
R_G_15_23_15_23  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_15_23_15_23  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA3-_Group_mid  4.507647e-20
R_G_15_24_15_24  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_15_24_15_24  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA4+_Group_mid  4.808995e-20
R_G_15_25_15_25  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_15_25_15_25  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA4-_Group_mid  4.843927e-20
R_G_15_26_15_26  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_15_26_15_26  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA5+_Group_mid  6.052163e-20
R_G_15_27_15_27  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_15_27_15_27  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA5-_Group_mid  5.800907e-20
R_G_15_28_15_28  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_15_28_15_28  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA6+_Group_mid  4.257044e-20
R_G_15_29_15_29  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_15_29_15_29  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA6-_Group_mid  4.398052e-20
R_G_15_30_15_30  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_15_30_15_30  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA7+_Group_mid  4.306822e-20
R_G_15_31_15_31  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_15_31_15_31  FCHIP_RXDATA7-_Group_mid FCHIP_TXDATA7-_Group_mid  4.412654e-20
C_16_17_16_17  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA0-_Group_mid  7.914042e-14
R_G_16_18_16_18  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA1+_Group_mid  2.841720e+08
C_16_18_16_18  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA1+_Group_mid  2.895033e-16
R_G_16_19_16_19  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA1-_Group_mid  1.000000e+09
C_16_19_16_19  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA1-_Group_mid  5.371526e-17
R_G_16_20_16_20  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_16_20_16_20  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA2+_Group_mid  9.116262e-19
R_G_16_21_16_21  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_16_21_16_21  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA2-_Group_mid  4.759955e-19
R_G_16_22_16_22  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_16_22_16_22  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA3+_Group_mid  8.182321e-20
R_G_16_23_16_23  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_16_23_16_23  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA3-_Group_mid  7.041022e-20
R_G_16_24_16_24  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_16_24_16_24  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA4+_Group_mid  7.763194e-20
R_G_16_25_16_25  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_16_25_16_25  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA4-_Group_mid  6.698131e-20
R_G_16_26_16_26  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_16_26_16_26  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA5+_Group_mid  7.287354e-20
R_G_16_27_16_27  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_16_27_16_27  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA5-_Group_mid  5.827932e-20
R_G_16_28_16_28  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_16_28_16_28  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA6+_Group_mid  4.963728e-20
R_G_16_29_16_29  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_16_29_16_29  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA6-_Group_mid  5.194067e-20
R_G_16_30_16_30  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_16_30_16_30  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA7+_Group_mid  5.165690e-20
R_G_16_31_16_31  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_16_31_16_31  FCHIP_TXDATA0+_Group_mid FCHIP_TXDATA7-_Group_mid  5.436115e-20
R_G_17_18_17_18  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA1+_Group_mid  9.317017e+07
C_17_18_17_18  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA1+_Group_mid  7.243260e-16
R_G_17_19_17_19  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA1-_Group_mid  3.021603e+08
C_17_19_17_19  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA1-_Group_mid  2.461838e-16
R_G_17_20_17_20  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA2+_Group_mid  1.000000e+09
C_17_20_17_20  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA2+_Group_mid  2.829806e-19
R_G_17_21_17_21  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA2-_Group_mid  1.000000e+09
C_17_21_17_21  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA2-_Group_mid  2.044231e-19
R_G_17_22_17_22  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_17_22_17_22  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA3+_Group_mid  2.358594e-19
R_G_17_23_17_23  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_17_23_17_23  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA3-_Group_mid  1.538939e-19
R_G_17_24_17_24  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_17_24_17_24  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA4+_Group_mid  1.852438e-19
R_G_17_25_17_25  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_17_25_17_25  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA4-_Group_mid  1.193213e-19
R_G_17_26_17_26  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_17_26_17_26  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA5+_Group_mid  1.899786e-19
R_G_17_27_17_27  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_17_27_17_27  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA5-_Group_mid  7.305579e-20
R_G_17_28_17_28  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_17_28_17_28  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA6+_Group_mid  4.878852e-20
R_G_17_29_17_29  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_17_29_17_29  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA6-_Group_mid  4.394376e-20
R_G_17_30_17_30  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_17_30_17_30  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA7+_Group_mid  4.910856e-20
R_G_17_31_17_31  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_17_31_17_31  FCHIP_TXDATA0-_Group_mid FCHIP_TXDATA7-_Group_mid  5.128406e-20
C_18_19_18_19  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA1-_Group_mid  9.096823e-14
R_G_18_20_18_20  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA2+_Group_mid  1.348362e+08
C_18_20_18_20  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA2+_Group_mid  4.834258e-16
R_G_18_21_18_21  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA2-_Group_mid  2.982727e+08
C_18_21_18_21  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA2-_Group_mid  2.512071e-16
R_G_18_22_18_22  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_18_22_18_22  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA3+_Group_mid  6.426358e-18
R_G_18_23_18_23  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_18_23_18_23  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA3-_Group_mid  1.547698e-17
R_G_18_24_18_24  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_18_24_18_24  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA4+_Group_mid  2.971373e-18
R_G_18_25_18_25  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_18_25_18_25  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA4-_Group_mid  1.585750e-19
R_G_18_26_18_26  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_18_26_18_26  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA5+_Group_mid  2.400894e-19
R_G_18_27_18_27  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_18_27_18_27  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA5-_Group_mid  1.709509e-18
R_G_18_28_18_28  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_18_28_18_28  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA6+_Group_mid  6.747271e-20
R_G_18_29_18_29  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_18_29_18_29  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA6-_Group_mid  4.390071e-20
R_G_18_30_18_30  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_18_30_18_30  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA7+_Group_mid  5.100833e-20
R_G_18_31_18_31  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_18_31_18_31  FCHIP_TXDATA1+_Group_mid FCHIP_TXDATA7-_Group_mid  5.739404e-20
R_G_19_20_19_20  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA2+_Group_mid  5.427394e+07
C_19_20_19_20  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA2+_Group_mid  1.155749e-15
R_G_19_21_19_21  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA2-_Group_mid  1.276736e+08
C_19_21_19_21  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA2-_Group_mid  5.367385e-16
R_G_19_22_19_22  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA3+_Group_mid  1.000000e+09
C_19_22_19_22  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA3+_Group_mid  1.215671e-17
R_G_19_23_19_23  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA3-_Group_mid  1.000000e+09
C_19_23_19_23  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA3-_Group_mid  2.760915e-17
R_G_19_24_19_24  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_19_24_19_24  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA4+_Group_mid  4.232759e-18
R_G_19_25_19_25  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_19_25_19_25  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA4-_Group_mid  2.225475e-19
R_G_19_26_19_26  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_19_26_19_26  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA5+_Group_mid  3.583241e-19
R_G_19_27_19_27  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_19_27_19_27  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA5-_Group_mid  1.999220e-18
R_G_19_28_19_28  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_19_28_19_28  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA6+_Group_mid  6.113643e-20
R_G_19_29_19_29  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_19_29_19_29  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA6-_Group_mid  5.726279e-20
R_G_19_30_19_30  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_19_30_19_30  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA7+_Group_mid  5.304199e-20
R_G_19_31_19_31  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_19_31_19_31  FCHIP_TXDATA1-_Group_mid FCHIP_TXDATA7-_Group_mid  5.989160e-20
C_20_21_20_21  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA2-_Group_mid  8.650563e-14
R_G_20_22_20_22  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA3+_Group_mid  1.875311e+08
C_20_22_20_22  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA3+_Group_mid  3.841886e-16
R_G_20_23_20_23  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA3-_Group_mid  3.507439e+08
C_20_23_20_23  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA3-_Group_mid  2.576630e-16
R_G_20_24_20_24  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_20_24_20_24  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA4+_Group_mid  1.670499e-17
R_G_20_25_20_25  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_20_25_20_25  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA4-_Group_mid  9.672728e-18
R_G_20_26_20_26  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_20_26_20_26  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA5+_Group_mid  9.778718e-19
R_G_20_27_20_27  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_20_27_20_27  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA5-_Group_mid  9.167355e-19
R_G_20_28_20_28  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_20_28_20_28  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA6+_Group_mid  5.577660e-20
R_G_20_29_20_29  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_20_29_20_29  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA6-_Group_mid  5.335621e-20
R_G_20_30_20_30  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_20_30_20_30  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA7+_Group_mid  4.748708e-20
R_G_20_31_20_31  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_20_31_20_31  FCHIP_TXDATA2+_Group_mid FCHIP_TXDATA7-_Group_mid  5.987221e-20
R_G_21_22_21_22  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA3+_Group_mid  6.596245e+07
C_21_22_21_22  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA3+_Group_mid  1.044025e-15
R_G_21_23_21_23  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA3-_Group_mid  9.295538e+07
C_21_23_21_23  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA3-_Group_mid  8.652175e-16
R_G_21_24_21_24  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA4+_Group_mid  1.000000e+09
C_21_24_21_24  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA4+_Group_mid  8.742579e-17
R_G_21_25_21_25  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA4-_Group_mid  1.000000e+09
C_21_25_21_25  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA4-_Group_mid  2.148988e-17
R_G_21_26_21_26  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_21_26_21_26  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA5+_Group_mid  1.738605e-18
R_G_21_27_21_27  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_21_27_21_27  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA5-_Group_mid  1.265560e-17
R_G_21_28_21_28  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_21_28_21_28  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA6+_Group_mid  7.484496e-20
R_G_21_29_21_29  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_21_29_21_29  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA6-_Group_mid  6.604759e-20
R_G_21_30_21_30  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_21_30_21_30  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA7+_Group_mid  6.141783e-20
R_G_21_31_21_31  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_21_31_21_31  FCHIP_TXDATA2-_Group_mid FCHIP_TXDATA7-_Group_mid  7.013576e-20
R_G_22_23_22_23  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA3-_Group_mid  1.079947e+06
C_22_23_22_23  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA3-_Group_mid  7.137031e-14
R_G_22_24_22_24  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA4+_Group_mid  6.689832e+07
C_22_24_22_24  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA4+_Group_mid  1.013956e-15
R_G_22_25_22_25  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA4-_Group_mid  1.824431e+08
C_22_25_22_25  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA4-_Group_mid  3.924730e-16
R_G_22_26_22_26  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_22_26_22_26  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA5+_Group_mid  1.273786e-17
R_G_22_27_22_27  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_22_27_22_27  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA5-_Group_mid  8.286760e-18
R_G_22_28_22_28  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_22_28_22_28  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA6+_Group_mid  5.498898e-20
R_G_22_29_22_29  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_22_29_22_29  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA6-_Group_mid  5.844708e-20
R_G_22_30_22_30  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_22_30_22_30  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA7+_Group_mid  4.918882e-20
R_G_22_31_22_31  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_22_31_22_31  FCHIP_TXDATA3+_Group_mid FCHIP_TXDATA7-_Group_mid  6.118324e-20
R_G_23_24_23_24  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA4+_Group_mid  1.782711e+07
C_23_24_23_24  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA4+_Group_mid  4.074434e-15
R_G_23_25_23_25  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA4-_Group_mid  6.211328e+07
C_23_25_23_25  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA4-_Group_mid  1.109177e-15
R_G_23_26_23_26  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA5+_Group_mid  1.000000e+09
C_23_26_23_26  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA5+_Group_mid  2.407469e-17
R_G_23_27_23_27  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA5-_Group_mid  1.000000e+09
C_23_27_23_27  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA5-_Group_mid  5.016169e-17
R_G_23_28_23_28  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_23_28_23_28  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA6+_Group_mid  8.899869e-20
R_G_23_29_23_29  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_23_29_23_29  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA6-_Group_mid  1.072832e-19
R_G_23_30_23_30  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_23_30_23_30  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA7+_Group_mid  5.411918e-20
R_G_23_31_23_31  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_23_31_23_31  FCHIP_TXDATA3-_Group_mid FCHIP_TXDATA7-_Group_mid  1.071999e-19
C_24_25_24_25  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA4-_Group_mid  1.043034e-13
R_G_24_26_24_26  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA5+_Group_mid  6.170960e+07
C_24_26_24_26  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA5+_Group_mid  1.146335e-15
R_G_24_27_24_27  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA5-_Group_mid  1.021294e+08
C_24_27_24_27  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA5-_Group_mid  7.875149e-16
R_G_24_28_24_28  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_24_28_24_28  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA6+_Group_mid  2.991829e-19
R_G_24_29_24_29  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_24_29_24_29  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA6-_Group_mid  2.141610e-19
R_G_24_30_24_30  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_24_30_24_30  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA7+_Group_mid  8.143345e-20
R_G_24_31_24_31  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_24_31_24_31  FCHIP_TXDATA4+_Group_mid FCHIP_TXDATA7-_Group_mid  1.662981e-19
R_G_25_26_25_26  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA5+_Group_mid  2.787814e+07
C_25_26_25_26  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA5+_Group_mid  2.394525e-15
R_G_25_27_25_27  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA5-_Group_mid  6.089711e+07
C_25_27_25_27  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA5-_Group_mid  1.160607e-15
R_G_25_28_25_28  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_25_28_25_28  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA6+_Group_mid  4.595354e-19
R_G_25_29_25_29  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_25_29_25_29  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA6-_Group_mid  3.189391e-19
R_G_25_30_25_30  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_25_30_25_30  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA7+_Group_mid  1.044521e-19
R_G_25_31_25_31  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_25_31_25_31  FCHIP_TXDATA4-_Group_mid FCHIP_TXDATA7-_Group_mid  2.510743e-19
C_26_27_26_27  FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA5-_Group_mid  1.162894e-13
R_G_26_28_26_28  FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_26_28_26_28  FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA6+_Group_mid  4.393757e-19
R_G_26_29_26_29  FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_26_29_26_29  FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA6-_Group_mid  7.932210e-19
R_G_26_30_26_30  FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_26_30_26_30  FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA7+_Group_mid  2.203218e-19
R_G_26_31_26_31  FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_26_31_26_31  FCHIP_TXDATA5+_Group_mid FCHIP_TXDATA7-_Group_mid  5.529545e-19
R_G_27_28_27_28  FCHIP_TXDATA5-_Group_mid FCHIP_TXDATA6+_Group_mid  1.000000e+09
C_27_28_27_28  FCHIP_TXDATA5-_Group_mid FCHIP_TXDATA6+_Group_mid  8.298549e-19
R_G_27_29_27_29  FCHIP_TXDATA5-_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_27_29_27_29  FCHIP_TXDATA5-_Group_mid FCHIP_TXDATA6-_Group_mid  1.232862e-18
R_G_27_30_27_30  FCHIP_TXDATA5-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_27_30_27_30  FCHIP_TXDATA5-_Group_mid FCHIP_TXDATA7+_Group_mid  4.792752e-19
R_G_27_31_27_31  FCHIP_TXDATA5-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_27_31_27_31  FCHIP_TXDATA5-_Group_mid FCHIP_TXDATA7-_Group_mid  8.128548e-19
R_G_28_29_28_29  FCHIP_TXDATA6+_Group_mid FCHIP_TXDATA6-_Group_mid  1.000000e+09
C_28_29_28_29  FCHIP_TXDATA6+_Group_mid FCHIP_TXDATA6-_Group_mid  1.304357e-18
R_G_28_30_28_30  FCHIP_TXDATA6+_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_28_30_28_30  FCHIP_TXDATA6+_Group_mid FCHIP_TXDATA7+_Group_mid  3.959102e-19
R_G_28_31_28_31  FCHIP_TXDATA6+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_28_31_28_31  FCHIP_TXDATA6+_Group_mid FCHIP_TXDATA7-_Group_mid  4.637228e-19
R_G_29_30_29_30  FCHIP_TXDATA6-_Group_mid FCHIP_TXDATA7+_Group_mid  1.000000e+09
C_29_30_29_30  FCHIP_TXDATA6-_Group_mid FCHIP_TXDATA7+_Group_mid  4.876437e-19
R_G_29_31_29_31  FCHIP_TXDATA6-_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_29_31_29_31  FCHIP_TXDATA6-_Group_mid FCHIP_TXDATA7-_Group_mid  6.854875e-19
R_G_30_31_30_31  FCHIP_TXDATA7+_Group_mid FCHIP_TXDATA7-_Group_mid  1.000000e+09
C_30_31_30_31  FCHIP_TXDATA7+_Group_mid FCHIP_TXDATA7-_Group_mid  3.735115e-19
.ends a0000_CPA_Sim_1
