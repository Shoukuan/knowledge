* contains one subcircuit for each unique part in design

.subckt COMP1_part 1 2
C1 1 2 1.000000e-08
.ends COMP1_part

