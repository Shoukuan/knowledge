* Path and file = D:\Persional\02 SIwave\07 CPA\Workflow\CPA Radhawk RLGC.siwaveresults\0000_CPA_Sim_1\0000_CPA_Sim_1_PDN_Channel\0000_CPA_Sim_1_CSP_BGA_BGA.sp

.subckt a0000_CPA_Sim_1_CSP_BGA_BGA
+ BGA_VSS_SINK_ BGA_VDD_15_SINK_
V1 BGA_VDD_15_SINK_ 0 1.500000e+00
V2 BGA_VSS_SINK_ 0 0.000000e+00
.ends a0000_CPA_Sim_1_CSP_BGA_BGA
