* Macro model for project = 0002_CPA_Sim_3

.subckt a0002_CPA_Sim_3
+ U2A5_GND_Group Group_602433-081_C2B2_GND_1 Group_602433-081_C3B10_GND_1
+ Group_A36096-108_C3L22_GND_1 Group_C83410-012_C3L15_GND_1
+ Group_C83410-012_C3L17_GND_1 Group_C83410-012_C3L18_GND_1
+ Group_C83410-012_C3L20_GND_1 Group_C83410-012_C3L24_GND_1
+ Group_C83410-012_C3L26_GND_1 Group_C83410-012_C3L28_GND_1
+ Group_C83410-012_C3L29_GND_1 Group_C97875-001_C3B11_GND_1
+ Group_C97875-001_C3B9_GND_1 Group_E16347-001_C2B12_GND_1
+ Group_E16347-001_C3B17_GND_1 U2A5_V1P0_S0_Group Group_602433-081_C2B2_V1P0_S0_2
+ Group_602433-081_C3B10_V1P0_S0_2 Group_A36096-108_C3L22_V1P0_S0_2
+ Group_C83410-012_C3L15_V1P0_S0_2 Group_C83410-012_C3L17_V1P0_S0_2
+ Group_C83410-012_C3L18_V1P0_S0_2 Group_C83410-012_C3L20_V1P0_S0_2
+ Group_C83410-012_C3L24_V1P0_S0_2 Group_C83410-012_C3L26_V1P0_S0_2
+ Group_C83410-012_C3L28_V1P0_S0_2 Group_C83410-012_C3L29_V1P0_S0_2
+ Group_C97875-001_C3B11_V1P0_S0_2 Group_C97875-001_C3B9_V1P0_S0_2
+ Group_E16347-001_C2B12_V1P0_S0_2 Group_E16347-001_C3B17_V1P0_S0_2
+ XW_V1P0_S0_SINK_ XW_GND_SINK_

L1_0_0 U2A5_GND_Group U2A5_GND_Group_mid 1.288378e-09
L2_0_0 U2A5_GND_Group_mid U2A5_GND_Group_resist 1.288378e-09
L1_1_1 Group_602433-081_C2B2_GND_1 Group_602433-081_C2B2_GND_1_mid 0.000000e+00
L2_1_1 Group_602433-081_C2B2_GND_1_mid Group_602433-081_C2B2_GND_1_resist 0.000000e+00
L1_2_2 Group_602433-081_C3B10_GND_1 Group_602433-081_C3B10_GND_1_mid 0.000000e+00
L2_2_2 Group_602433-081_C3B10_GND_1_mid Group_602433-081_C3B10_GND_1_resist 0.000000e+00
L1_3_3 Group_A36096-108_C3L22_GND_1 Group_A36096-108_C3L22_GND_1_mid 0.000000e+00
L2_3_3 Group_A36096-108_C3L22_GND_1_mid Group_A36096-108_C3L22_GND_1_resist 0.000000e+00
L1_4_4 Group_C83410-012_C3L15_GND_1 Group_C83410-012_C3L15_GND_1_mid 0.000000e+00
L2_4_4 Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L15_GND_1_resist 0.000000e+00
L1_5_5 Group_C83410-012_C3L17_GND_1 Group_C83410-012_C3L17_GND_1_mid 0.000000e+00
L2_5_5 Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L17_GND_1_resist 0.000000e+00
L1_6_6 Group_C83410-012_C3L18_GND_1 Group_C83410-012_C3L18_GND_1_mid 0.000000e+00
L2_6_6 Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L18_GND_1_resist 0.000000e+00
L1_7_7 Group_C83410-012_C3L20_GND_1 Group_C83410-012_C3L20_GND_1_mid 0.000000e+00
L2_7_7 Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L20_GND_1_resist 0.000000e+00
L1_8_8 Group_C83410-012_C3L24_GND_1 Group_C83410-012_C3L24_GND_1_mid 0.000000e+00
L2_8_8 Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L24_GND_1_resist 0.000000e+00
L1_9_9 Group_C83410-012_C3L26_GND_1 Group_C83410-012_C3L26_GND_1_mid 0.000000e+00
L2_9_9 Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L26_GND_1_resist 0.000000e+00
L1_10_10 Group_C83410-012_C3L28_GND_1 Group_C83410-012_C3L28_GND_1_mid 0.000000e+00
L2_10_10 Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L28_GND_1_resist 0.000000e+00
L1_11_11 Group_C83410-012_C3L29_GND_1 Group_C83410-012_C3L29_GND_1_mid 0.000000e+00
L2_11_11 Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L29_GND_1_resist 0.000000e+00
L1_12_12 Group_C97875-001_C3B11_GND_1 Group_C97875-001_C3B11_GND_1_mid 0.000000e+00
L2_12_12 Group_C97875-001_C3B11_GND_1_mid Group_C97875-001_C3B11_GND_1_resist 0.000000e+00
L1_13_13 Group_C97875-001_C3B9_GND_1 Group_C97875-001_C3B9_GND_1_mid 0.000000e+00
L2_13_13 Group_C97875-001_C3B9_GND_1_mid Group_C97875-001_C3B9_GND_1_resist 0.000000e+00
L1_14_14 Group_E16347-001_C2B12_GND_1 Group_E16347-001_C2B12_GND_1_mid 0.000000e+00
L2_14_14 Group_E16347-001_C2B12_GND_1_mid Group_E16347-001_C2B12_GND_1_resist 0.000000e+00
L1_15_15 Group_E16347-001_C3B17_GND_1 Group_E16347-001_C3B17_GND_1_mid 0.000000e+00
L2_15_15 Group_E16347-001_C3B17_GND_1_mid Group_E16347-001_C3B17_GND_1_resist 0.000000e+00
L1_16_16 U2A5_V1P0_S0_Group U2A5_V1P0_S0_Group_mid 1.317516e-09
L2_16_16 U2A5_V1P0_S0_Group_mid U2A5_V1P0_S0_Group_resist 1.317516e-09
L1_17_17 Group_602433-081_C2B2_V1P0_S0_2 Group_602433-081_C2B2_V1P0_S0_2_mid 9.647277e-10
L2_17_17 Group_602433-081_C2B2_V1P0_S0_2_mid Group_602433-081_C2B2_V1P0_S0_2_resist 9.647277e-10
L1_18_18 Group_602433-081_C3B10_V1P0_S0_2 Group_602433-081_C3B10_V1P0_S0_2_mid 3.680217e-10
L2_18_18 Group_602433-081_C3B10_V1P0_S0_2_mid Group_602433-081_C3B10_V1P0_S0_2_resist 3.680217e-10
L1_19_19 Group_A36096-108_C3L22_V1P0_S0_2 Group_A36096-108_C3L22_V1P0_S0_2_mid 1.406912e-09
L2_19_19 Group_A36096-108_C3L22_V1P0_S0_2_mid Group_A36096-108_C3L22_V1P0_S0_2_resist 1.406912e-09
L1_20_20 Group_C83410-012_C3L15_V1P0_S0_2 Group_C83410-012_C3L15_V1P0_S0_2_mid 1.170971e-09
L2_20_20 Group_C83410-012_C3L15_V1P0_S0_2_mid Group_C83410-012_C3L15_V1P0_S0_2_resist 1.170971e-09
L1_21_21 Group_C83410-012_C3L17_V1P0_S0_2 Group_C83410-012_C3L17_V1P0_S0_2_mid 1.315769e-09
L2_21_21 Group_C83410-012_C3L17_V1P0_S0_2_mid Group_C83410-012_C3L17_V1P0_S0_2_resist 1.315769e-09
L1_22_22 Group_C83410-012_C3L18_V1P0_S0_2 Group_C83410-012_C3L18_V1P0_S0_2_mid 1.356556e-09
L2_22_22 Group_C83410-012_C3L18_V1P0_S0_2_mid Group_C83410-012_C3L18_V1P0_S0_2_resist 1.356556e-09
L1_23_23 Group_C83410-012_C3L20_V1P0_S0_2 Group_C83410-012_C3L20_V1P0_S0_2_mid 1.341875e-09
L2_23_23 Group_C83410-012_C3L20_V1P0_S0_2_mid Group_C83410-012_C3L20_V1P0_S0_2_resist 1.341875e-09
L1_24_24 Group_C83410-012_C3L24_V1P0_S0_2 Group_C83410-012_C3L24_V1P0_S0_2_mid 1.324130e-09
L2_24_24 Group_C83410-012_C3L24_V1P0_S0_2_mid Group_C83410-012_C3L24_V1P0_S0_2_resist 1.324130e-09
L1_25_25 Group_C83410-012_C3L26_V1P0_S0_2 Group_C83410-012_C3L26_V1P0_S0_2_mid 1.309709e-09
L2_25_25 Group_C83410-012_C3L26_V1P0_S0_2_mid Group_C83410-012_C3L26_V1P0_S0_2_resist 1.309709e-09
L1_26_26 Group_C83410-012_C3L28_V1P0_S0_2 Group_C83410-012_C3L28_V1P0_S0_2_mid 1.343730e-09
L2_26_26 Group_C83410-012_C3L28_V1P0_S0_2_mid Group_C83410-012_C3L28_V1P0_S0_2_resist 1.343730e-09
L1_27_27 Group_C83410-012_C3L29_V1P0_S0_2 Group_C83410-012_C3L29_V1P0_S0_2_mid 1.335471e-09
L2_27_27 Group_C83410-012_C3L29_V1P0_S0_2_mid Group_C83410-012_C3L29_V1P0_S0_2_resist 1.335471e-09
L1_28_28 Group_C97875-001_C3B11_V1P0_S0_2 Group_C97875-001_C3B11_V1P0_S0_2_mid 1.326572e-09
L2_28_28 Group_C97875-001_C3B11_V1P0_S0_2_mid Group_C97875-001_C3B11_V1P0_S0_2_resist 1.326572e-09
L1_29_29 Group_C97875-001_C3B9_V1P0_S0_2 Group_C97875-001_C3B9_V1P0_S0_2_mid 1.337589e-09
L2_29_29 Group_C97875-001_C3B9_V1P0_S0_2_mid Group_C97875-001_C3B9_V1P0_S0_2_resist 1.337589e-09
L1_30_30 Group_E16347-001_C2B12_V1P0_S0_2 Group_E16347-001_C2B12_V1P0_S0_2_mid 6.763435e-10
L2_30_30 Group_E16347-001_C2B12_V1P0_S0_2_mid Group_E16347-001_C2B12_V1P0_S0_2_resist 6.763435e-10
L1_31_31 Group_E16347-001_C3B17_V1P0_S0_2 Group_E16347-001_C3B17_V1P0_S0_2_mid 6.625706e-10
L2_31_31 Group_E16347-001_C3B17_V1P0_S0_2_mid Group_E16347-001_C3B17_V1P0_S0_2_resist 6.625706e-10


R_d_1 Group_602433-081_C2B2_GND_1_resist Group_602433-081_C3B10_GND_1_resist 3.129651e-02
R_d_2 Group_602433-081_C2B2_GND_1_resist Group_A36096-108_C3L22_GND_1_resist 6.162747e-01
R_d_3 Group_602433-081_C2B2_GND_1_resist Group_C83410-012_C3L15_GND_1_resist 2.018983e+00
R_d_4 Group_602433-081_C2B2_GND_1_resist Group_C83410-012_C3L17_GND_1_resist 3.415827e+00
R_d_5 Group_602433-081_C2B2_GND_1_resist Group_C83410-012_C3L18_GND_1_resist 1.566836e+00
R_d_6 Group_602433-081_C2B2_GND_1_resist Group_C83410-012_C3L20_GND_1_resist 1.127169e+00
R_d_7 Group_602433-081_C2B2_GND_1_resist Group_C83410-012_C3L24_GND_1_resist 6.559219e-01
R_d_8 Group_602433-081_C2B2_GND_1_resist Group_C83410-012_C3L26_GND_1_resist 5.257978e-01
R_d_9 Group_602433-081_C2B2_GND_1_resist Group_C83410-012_C3L28_GND_1_resist 2.932697e-01
R_d_10 Group_602433-081_C2B2_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 4.173766e-01
R_d_11 Group_602433-081_C2B2_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 2.978453e-02
R_d_12 Group_602433-081_C2B2_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 3.106918e-02
R_d_13 Group_602433-081_C2B2_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 9.888440e-03
R_d_14 Group_602433-081_C2B2_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 5.697217e-02
R_d_15 Group_602433-081_C2B2_GND_1_resist XW_GND_SINK_ 3.641617e-02
R_d_16 Group_602433-081_C2B2_V1P0_S0_2_resist Group_602433-081_C3B10_V1P0_S0_2_resist 1.171072e-02
R_d_17 Group_602433-081_C2B2_V1P0_S0_2_resist Group_A36096-108_C3L22_V1P0_S0_2_resist 5.273684e-01
R_d_18 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C83410-012_C3L15_V1P0_S0_2_resist 1.375314e+00
R_d_19 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C83410-012_C3L17_V1P0_S0_2_resist 9.812274e-01
R_d_20 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C83410-012_C3L18_V1P0_S0_2_resist 2.048753e-01
R_d_21 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C83410-012_C3L20_V1P0_S0_2_resist 5.398154e-01
R_d_22 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C83410-012_C3L24_V1P0_S0_2_resist 1.611058e-01
R_d_23 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C83410-012_C3L26_V1P0_S0_2_resist 6.761194e-01
R_d_24 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 1.954631e-01
R_d_25 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 2.105836e-01
R_d_26 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 2.284273e-02
R_d_27 Group_602433-081_C2B2_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 1.730341e-02
R_d_28 Group_602433-081_C2B2_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 2.296554e-03
R_d_29 Group_602433-081_C2B2_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 9.118348e-03
R_d_30 Group_602433-081_C2B2_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 4.283272e-02
R_d_31 Group_602433-081_C3B10_GND_1_resist Group_A36096-108_C3L22_GND_1_resist 1.347596e+00
R_d_32 Group_602433-081_C3B10_GND_1_resist Group_C83410-012_C3L15_GND_1_resist 2.429429e+00
R_d_33 Group_602433-081_C3B10_GND_1_resist Group_C83410-012_C3L17_GND_1_resist 4.230324e+00
R_d_34 Group_602433-081_C3B10_GND_1_resist Group_C83410-012_C3L18_GND_1_resist 1.330560e+00
R_d_35 Group_602433-081_C3B10_GND_1_resist Group_C83410-012_C3L20_GND_1_resist 1.481044e+00
R_d_36 Group_602433-081_C3B10_GND_1_resist Group_C83410-012_C3L24_GND_1_resist 8.308564e-01
R_d_37 Group_602433-081_C3B10_GND_1_resist Group_C83410-012_C3L26_GND_1_resist 1.080668e+00
R_d_38 Group_602433-081_C3B10_GND_1_resist Group_C83410-012_C3L28_GND_1_resist 4.259490e-01
R_d_39 Group_602433-081_C3B10_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 6.919924e-01
R_d_40 Group_602433-081_C3B10_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 1.899076e-02
R_d_41 Group_602433-081_C3B10_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 1.894571e-02
R_d_42 Group_602433-081_C3B10_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 1.575309e-02
R_d_43 Group_602433-081_C3B10_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 2.909375e-02
R_d_44 Group_602433-081_C3B10_GND_1_resist XW_GND_SINK_ 2.472492e-02
R_d_45 Group_602433-081_C3B10_V1P0_S0_2_resist Group_A36096-108_C3L22_V1P0_S0_2_resist 8.896194e-01
R_d_46 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C83410-012_C3L15_V1P0_S0_2_resist 2.312435e+00
R_d_47 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C83410-012_C3L17_V1P0_S0_2_resist 1.650995e+00
R_d_48 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C83410-012_C3L18_V1P0_S0_2_resist 3.446324e-01
R_d_49 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C83410-012_C3L20_V1P0_S0_2_resist 9.081936e-01
R_d_50 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C83410-012_C3L24_V1P0_S0_2_resist 2.712154e-01
R_d_51 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C83410-012_C3L26_V1P0_S0_2_resist 1.141981e+00
R_d_52 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 3.303456e-01
R_d_53 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 3.560144e-01
R_d_54 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 1.049102e-02
R_d_55 Group_602433-081_C3B10_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 7.885120e-03
R_d_56 Group_602433-081_C3B10_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 1.152338e-02
R_d_57 Group_602433-081_C3B10_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 1.257997e-02
R_d_58 Group_602433-081_C3B10_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 1.984497e-02
R_d_59 Group_A36096-108_C3L22_GND_1_resist Group_C83410-012_C3L15_GND_1_resist 2.391814e-02
R_d_60 Group_A36096-108_C3L22_GND_1_resist Group_C83410-012_C3L17_GND_1_resist 3.797684e-02
R_d_61 Group_A36096-108_C3L22_GND_1_resist Group_C83410-012_C3L18_GND_1_resist 1.191512e-01
R_d_62 Group_A36096-108_C3L22_GND_1_resist Group_C83410-012_C3L20_GND_1_resist 2.938456e-02
R_d_63 Group_A36096-108_C3L22_GND_1_resist Group_C83410-012_C3L24_GND_1_resist 9.859195e-02
R_d_64 Group_A36096-108_C3L22_GND_1_resist Group_C83410-012_C3L26_GND_1_resist 2.320009e-03
R_d_65 Group_A36096-108_C3L22_GND_1_resist Group_C83410-012_C3L28_GND_1_resist 4.293529e-02
R_d_66 Group_A36096-108_C3L22_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 9.546949e-03
R_d_67 Group_A36096-108_C3L22_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 1.191854e+00
R_d_68 Group_A36096-108_C3L22_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 1.254447e+00
R_d_69 Group_A36096-108_C3L22_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 4.987157e-01
R_d_70 Group_A36096-108_C3L22_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 1.376878e+00
R_d_71 Group_A36096-108_C3L22_GND_1_resist XW_GND_SINK_ 1.398339e+00
R_d_72 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C83410-012_C3L15_V1P0_S0_2_resist 1.082866e-02
R_d_73 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C83410-012_C3L17_V1P0_S0_2_resist 2.763793e-03
R_d_74 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C83410-012_C3L18_V1P0_S0_2_resist 1.112869e-02
R_d_75 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C83410-012_C3L20_V1P0_S0_2_resist 2.246385e-03
R_d_76 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C83410-012_C3L24_V1P0_S0_2_resist 2.472210e-02
R_d_77 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C83410-012_C3L26_V1P0_S0_2_resist 1.171591e-03
R_d_78 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 9.413553e-03
R_d_79 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 7.780664e-03
R_d_80 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 1.829197e+00
R_d_81 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 1.382788e+00
R_d_82 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 5.001081e-01
R_d_83 Group_A36096-108_C3L22_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 2.598723e-01
R_d_84 Group_A36096-108_C3L22_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 3.437763e+00
R_d_85 Group_C83410-012_C3L15_GND_1_resist Group_C83410-012_C3L17_GND_1_resist 1.056767e-03
R_d_86 Group_C83410-012_C3L15_GND_1_resist Group_C83410-012_C3L18_GND_1_resist 1.567104e-02
R_d_87 Group_C83410-012_C3L15_GND_1_resist Group_C83410-012_C3L20_GND_1_resist 5.339605e-02
R_d_88 Group_C83410-012_C3L15_GND_1_resist Group_C83410-012_C3L24_GND_1_resist 2.150921e-01
R_d_89 Group_C83410-012_C3L15_GND_1_resist Group_C83410-012_C3L26_GND_1_resist 7.256187e-02
R_d_90 Group_C83410-012_C3L15_GND_1_resist Group_C83410-012_C3L28_GND_1_resist 1.982852e-01
R_d_91 Group_C83410-012_C3L15_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 1.696813e-01
R_d_92 Group_C83410-012_C3L15_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 8.538087e-01
R_d_93 Group_C83410-012_C3L15_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 9.674166e-01
R_d_94 Group_C83410-012_C3L15_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 1.457560e+00
R_d_95 Group_C83410-012_C3L15_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 1.577613e+00
R_d_96 Group_C83410-012_C3L15_GND_1_resist XW_GND_SINK_ 8.597921e-01
R_d_97 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_C83410-012_C3L17_V1P0_S0_2_resist 6.250385e-03
R_d_98 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_C83410-012_C3L18_V1P0_S0_2_resist 1.304318e-02
R_d_99 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_C83410-012_C3L20_V1P0_S0_2_resist 3.857695e-03
R_d_100 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_C83410-012_C3L24_V1P0_S0_2_resist 6.803984e-02
R_d_101 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_C83410-012_C3L26_V1P0_S0_2_resist 6.202149e-02
R_d_102 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 1.611991e-01
R_d_103 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 1.730848e-01
R_d_104 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 4.755738e+00
R_d_105 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 3.595085e+00
R_d_106 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 1.304345e+00
R_d_107 Group_C83410-012_C3L15_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 6.691899e-01
R_d_108 Group_C83410-012_C3L15_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 8.937948e+00
R_d_109 Group_C83410-012_C3L17_GND_1_resist Group_C83410-012_C3L18_GND_1_resist 2.735495e-02
R_d_110 Group_C83410-012_C3L17_GND_1_resist Group_C83410-012_C3L20_GND_1_resist 9.205215e-02
R_d_111 Group_C83410-012_C3L17_GND_1_resist Group_C83410-012_C3L24_GND_1_resist 3.768068e-01
R_d_112 Group_C83410-012_C3L17_GND_1_resist Group_C83410-012_C3L26_GND_1_resist 1.164201e-01
R_d_113 Group_C83410-012_C3L17_GND_1_resist Group_C83410-012_C3L28_GND_1_resist 3.439355e-01
R_d_114 Group_C83410-012_C3L17_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 2.804481e-01
R_d_115 Group_C83410-012_C3L17_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 1.508100e+00
R_d_116 Group_C83410-012_C3L17_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 1.708087e+00
R_d_117 Group_C83410-012_C3L17_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 2.489379e+00
R_d_118 Group_C83410-012_C3L17_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 2.782943e+00
R_d_119 Group_C83410-012_C3L17_GND_1_resist XW_GND_SINK_ 1.519733e+00
R_d_120 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_C83410-012_C3L18_V1P0_S0_2_resist 1.319304e-02
R_d_121 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_C83410-012_C3L20_V1P0_S0_2_resist 3.085439e-03
R_d_122 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_C83410-012_C3L24_V1P0_S0_2_resist 5.241561e-02
R_d_123 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_C83410-012_C3L26_V1P0_S0_2_resist 1.766504e-02
R_d_124 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 7.601361e-02
R_d_125 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 7.364202e-02
R_d_126 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 3.395270e+00
R_d_127 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 2.566648e+00
R_d_128 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 9.305752e-01
R_d_129 Group_C83410-012_C3L17_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 4.787462e-01
R_d_130 Group_C83410-012_C3L17_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 6.381066e+00
R_d_131 Group_C83410-012_C3L18_GND_1_resist Group_C83410-012_C3L20_GND_1_resist 8.334412e-03
R_d_132 Group_C83410-012_C3L18_GND_1_resist Group_C83410-012_C3L24_GND_1_resist 3.920386e-02
R_d_133 Group_C83410-012_C3L18_GND_1_resist Group_C83410-012_C3L26_GND_1_resist 1.004405e-01
R_d_134 Group_C83410-012_C3L18_GND_1_resist Group_C83410-012_C3L28_GND_1_resist 4.069892e-02
R_d_135 Group_C83410-012_C3L18_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 6.594089e-02
R_d_136 Group_C83410-012_C3L18_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 5.252359e-01
R_d_137 Group_C83410-012_C3L18_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 5.770707e-01
R_d_138 Group_C83410-012_C3L18_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 9.415369e-01
R_d_139 Group_C83410-012_C3L18_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 6.926516e-01
R_d_140 Group_C83410-012_C3L18_GND_1_resist XW_GND_SINK_ 5.626392e-01
R_d_141 Group_C83410-012_C3L18_V1P0_S0_2_resist Group_C83410-012_C3L20_V1P0_S0_2_resist 1.108942e-03
R_d_142 Group_C83410-012_C3L18_V1P0_S0_2_resist Group_C83410-012_C3L24_V1P0_S0_2_resist 2.382705e-03
R_d_143 Group_C83410-012_C3L18_V1P0_S0_2_resist Group_C83410-012_C3L26_V1P0_S0_2_resist 3.721481e-02
R_d_144 Group_C83410-012_C3L18_V1P0_S0_2_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 1.228970e-02
R_d_145 Group_C83410-012_C3L18_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 1.699002e-02
R_d_146 Group_C83410-012_C3L18_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 7.087477e-01
R_d_147 Group_C83410-012_C3L18_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 5.357762e-01
R_d_148 Group_C83410-012_C3L18_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 1.943008e-01
R_d_149 Group_C83410-012_C3L18_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 9.986281e-02
R_d_150 Group_C83410-012_C3L18_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 1.332021e+00
R_d_151 Group_C83410-012_C3L20_GND_1_resist Group_C83410-012_C3L24_GND_1_resist 1.075513e-02
R_d_152 Group_C83410-012_C3L20_GND_1_resist Group_C83410-012_C3L26_GND_1_resist 1.394274e-02
R_d_153 Group_C83410-012_C3L20_GND_1_resist Group_C83410-012_C3L28_GND_1_resist 1.097229e-02
R_d_154 Group_C83410-012_C3L20_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 1.040818e-02
R_d_155 Group_C83410-012_C3L20_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 8.818568e-01
R_d_156 Group_C83410-012_C3L20_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 9.434310e-01
R_d_157 Group_C83410-012_C3L20_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 7.571160e-01
R_d_158 Group_C83410-012_C3L20_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 9.523319e-01
R_d_159 Group_C83410-012_C3L20_GND_1_resist XW_GND_SINK_ 9.974379e-01
R_d_160 Group_C83410-012_C3L20_V1P0_S0_2_resist Group_C83410-012_C3L24_V1P0_S0_2_resist 8.909159e-03
R_d_161 Group_C83410-012_C3L20_V1P0_S0_2_resist Group_C83410-012_C3L26_V1P0_S0_2_resist 1.505621e-02
R_d_162 Group_C83410-012_C3L20_V1P0_S0_2_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 3.147946e-02
R_d_163 Group_C83410-012_C3L20_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 3.681672e-02
R_d_164 Group_C83410-012_C3L20_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 1.867711e+00
R_d_165 Group_C83410-012_C3L20_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 1.411892e+00
R_d_166 Group_C83410-012_C3L20_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 5.119510e-01
R_d_167 Group_C83410-012_C3L20_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 2.632786e-01
R_d_168 Group_C83410-012_C3L20_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 3.510175e+00
R_d_169 Group_C83410-012_C3L24_GND_1_resist Group_C83410-012_C3L26_GND_1_resist 4.620357e-02
R_d_170 Group_C83410-012_C3L24_GND_1_resist Group_C83410-012_C3L28_GND_1_resist 1.830564e-03
R_d_171 Group_C83410-012_C3L24_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 1.163422e-02
R_d_172 Group_C83410-012_C3L24_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 5.307061e-01
R_d_173 Group_C83410-012_C3L24_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 5.624077e-01
R_d_174 Group_C83410-012_C3L24_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 4.271894e-01
R_d_175 Group_C83410-012_C3L24_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 5.228116e-01
R_d_176 Group_C83410-012_C3L24_GND_1_resist XW_GND_SINK_ 6.126069e-01
R_d_177 Group_C83410-012_C3L24_V1P0_S0_2_resist Group_C83410-012_C3L26_V1P0_S0_2_resist 3.154956e-02
R_d_178 Group_C83410-012_C3L24_V1P0_S0_2_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 5.541738e-03
R_d_179 Group_C83410-012_C3L24_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 7.989652e-03
R_d_180 Group_C83410-012_C3L24_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 5.577352e-01
R_d_181 Group_C83410-012_C3L24_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 4.216196e-01
R_d_182 Group_C83410-012_C3L24_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 1.527870e-01
R_d_183 Group_C83410-012_C3L24_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 7.876334e-02
R_d_184 Group_C83410-012_C3L24_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 1.048205e+00
R_d_185 Group_C83410-012_C3L26_GND_1_resist Group_C83410-012_C3L28_GND_1_resist 1.932686e-02
R_d_186 Group_C83410-012_C3L26_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 1.915102e-03
R_d_187 Group_C83410-012_C3L26_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 9.927528e-01
R_d_188 Group_C83410-012_C3L26_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 1.035694e+00
R_d_189 Group_C83410-012_C3L26_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 4.109210e-01
R_d_190 Group_C83410-012_C3L26_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 1.045325e+00
R_d_191 Group_C83410-012_C3L26_GND_1_resist XW_GND_SINK_ 1.188515e+00
R_d_192 Group_C83410-012_C3L26_V1P0_S0_2_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 8.238032e-03
R_d_193 Group_C83410-012_C3L26_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 6.678678e-03
R_d_194 Group_C83410-012_C3L26_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 2.347901e+00
R_d_195 Group_C83410-012_C3L26_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 1.774911e+00
R_d_196 Group_C83410-012_C3L26_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 6.411468e-01
R_d_197 Group_C83410-012_C3L26_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 3.348044e-01
R_d_198 Group_C83410-012_C3L26_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 4.412589e+00
R_d_199 Group_C83410-012_C3L28_GND_1_resist Group_C83410-012_C3L29_GND_1_resist 3.160042e-03
R_d_200 Group_C83410-012_C3L28_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 3.233825e-01
R_d_201 Group_C83410-012_C3L28_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 3.391886e-01
R_d_202 Group_C83410-012_C3L28_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 1.974105e-01
R_d_203 Group_C83410-012_C3L28_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 3.045611e-01
R_d_204 Group_C83410-012_C3L28_GND_1_resist XW_GND_SINK_ 3.817684e-01
R_d_205 Group_C83410-012_C3L28_V1P0_S0_2_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 9.794370e-04
R_d_206 Group_C83410-012_C3L28_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 6.791598e-01
R_d_207 Group_C83410-012_C3L28_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 5.134161e-01
R_d_208 Group_C83410-012_C3L28_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 1.853494e-01
R_d_209 Group_C83410-012_C3L28_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 9.702400e-02
R_d_210 Group_C83410-012_C3L28_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 1.276394e+00
R_d_211 Group_C83410-012_C3L29_GND_1_resist Group_C97875-001_C3B11_GND_1_resist 5.819444e-01
R_d_212 Group_C83410-012_C3L29_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 6.073832e-01
R_d_213 Group_C83410-012_C3L29_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 2.955879e-01
R_d_214 Group_C83410-012_C3L29_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 5.552544e-01
R_d_215 Group_C83410-012_C3L29_GND_1_resist XW_GND_SINK_ 6.950099e-01
R_d_216 Group_C83410-012_C3L29_V1P0_S0_2_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 7.319172e-01
R_d_217 Group_C83410-012_C3L29_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 5.532989e-01
R_d_218 Group_C83410-012_C3L29_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 1.996857e-01
R_d_219 Group_C83410-012_C3L29_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 1.046605e-01
R_d_220 Group_C83410-012_C3L29_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 1.375544e+00
R_d_221 Group_C97875-001_C3B11_GND_1_resist Group_C97875-001_C3B9_GND_1_resist 7.487758e-04
R_d_222 Group_C97875-001_C3B11_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 1.841842e-02
R_d_223 Group_C97875-001_C3B11_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 2.431993e-02
R_d_224 Group_C97875-001_C3B11_GND_1_resist XW_GND_SINK_ 2.945246e-03
R_d_225 Group_C97875-001_C3B11_V1P0_S0_2_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 6.416349e-04
R_d_226 Group_C97875-001_C3B11_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 2.256395e-02
R_d_227 Group_C97875-001_C3B11_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 2.620051e-02
R_d_228 Group_C97875-001_C3B11_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 1.270723e-03
R_d_229 Group_C97875-001_C3B9_GND_1_resist Group_E16347-001_C2B12_GND_1_resist 1.893497e-02
R_d_230 Group_C97875-001_C3B9_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 2.429532e-02
R_d_231 Group_C97875-001_C3B9_GND_1_resist XW_GND_SINK_ 4.337281e-03
R_d_232 Group_C97875-001_C3B9_V1P0_S0_2_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 1.708992e-02
R_d_233 Group_C97875-001_C3B9_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 1.979508e-02
R_d_234 Group_C97875-001_C3B9_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 2.169785e-03
R_d_235 Group_E16347-001_C2B12_GND_1_resist Group_E16347-001_C3B17_GND_1_resist 2.792484e-02
R_d_236 Group_E16347-001_C2B12_GND_1_resist XW_GND_SINK_ 2.297823e-02
R_d_237 Group_E16347-001_C2B12_V1P0_S0_2_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 8.701845e-03
R_d_238 Group_E16347-001_C2B12_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 4.231636e-02
R_d_239 Group_E16347-001_C3B17_GND_1_resist XW_GND_SINK_ 3.151707e-02
R_d_240 Group_E16347-001_C3B17_V1P0_S0_2_resist XW_V1P0_S0_SINK_ 4.927205e-02
R_d_241 U2A5_GND_Group_resist Group_602433-081_C2B2_GND_1_resist 3.528042e-03
R_d_242 U2A5_GND_Group_resist Group_602433-081_C3B10_GND_1_resist 4.149212e-03
R_d_243 U2A5_GND_Group_resist Group_A36096-108_C3L22_GND_1_resist 4.416357e-04
R_d_244 U2A5_GND_Group_resist Group_C83410-012_C3L15_GND_1_resist 6.025860e-04
R_d_245 U2A5_GND_Group_resist Group_C83410-012_C3L17_GND_1_resist 1.022445e-03
R_d_246 U2A5_GND_Group_resist Group_C83410-012_C3L18_GND_1_resist 7.673083e-04
R_d_247 U2A5_GND_Group_resist Group_C83410-012_C3L20_GND_1_resist 1.404689e-03
R_d_248 U2A5_GND_Group_resist Group_C83410-012_C3L24_GND_1_resist 1.072334e-03
R_d_249 U2A5_GND_Group_resist Group_C83410-012_C3L26_GND_1_resist 6.179431e-04
R_d_250 U2A5_GND_Group_resist Group_C83410-012_C3L28_GND_1_resist 6.503350e-04
R_d_251 U2A5_GND_Group_resist Group_C83410-012_C3L29_GND_1_resist 7.625357e-04
R_d_252 U2A5_GND_Group_resist Group_C97875-001_C3B11_GND_1_resist 2.287160e-03
R_d_253 U2A5_GND_Group_resist Group_C97875-001_C3B9_GND_1_resist 2.480282e-03
R_d_254 U2A5_GND_Group_resist Group_E16347-001_C2B12_GND_1_resist 2.303765e-03
R_d_255 U2A5_GND_Group_resist Group_E16347-001_C3B17_GND_1_resist 2.411443e-03
R_d_256 U2A5_GND_Group_resist XW_GND_SINK_ 2.507419e-03
R_d_257 U2A5_V1P0_S0_Group_resist Group_602433-081_C2B2_V1P0_S0_2_resist 1.692570e-02
R_d_258 U2A5_V1P0_S0_Group_resist Group_602433-081_C3B10_V1P0_S0_2_resist 2.851731e-02
R_d_259 U2A5_V1P0_S0_Group_resist Group_A36096-108_C3L22_V1P0_S0_2_resist 6.559298e-04
R_d_260 U2A5_V1P0_S0_Group_resist Group_C83410-012_C3L15_V1P0_S0_2_resist 1.560854e-03
R_d_261 U2A5_V1P0_S0_Group_resist Group_C83410-012_C3L17_V1P0_S0_2_resist 6.352764e-04
R_d_262 U2A5_V1P0_S0_Group_resist Group_C83410-012_C3L18_V1P0_S0_2_resist 9.533963e-04
R_d_263 U2A5_V1P0_S0_Group_resist Group_C83410-012_C3L20_V1P0_S0_2_resist 9.498352e-04
R_d_264 U2A5_V1P0_S0_Group_resist Group_C83410-012_C3L24_V1P0_S0_2_resist 1.027034e-03
R_d_265 U2A5_V1P0_S0_Group_resist Group_C83410-012_C3L26_V1P0_S0_2_resist 1.157495e-03
R_d_266 U2A5_V1P0_S0_Group_resist Group_C83410-012_C3L28_V1P0_S0_2_resist 1.363325e-03
R_d_267 U2A5_V1P0_S0_Group_resist Group_C83410-012_C3L29_V1P0_S0_2_resist 1.444487e-03
R_d_268 U2A5_V1P0_S0_Group_resist Group_C97875-001_C3B11_V1P0_S0_2_resist 5.864068e-02
R_d_269 U2A5_V1P0_S0_Group_resist Group_C97875-001_C3B9_V1P0_S0_2_resist 4.432949e-02
R_d_270 U2A5_V1P0_S0_Group_resist Group_E16347-001_C2B12_V1P0_S0_2_resist 1.605135e-02
R_d_271 U2A5_V1P0_S0_Group_resist Group_E16347-001_C3B17_V1P0_S0_2_resist 8.301280e-03
R_d_272 U2A5_V1P0_S0_Group_resist XW_V1P0_S0_SINK_ 1.102088e-01
K1_0_16  L1_0_0  L1_16_16  7.113024e-01
K2_0_16  L2_0_0  L2_16_16  7.113024e-01
K1_0_17  L1_0_0  L1_17_17  -7.218785e-01
K2_0_17  L2_0_0  L2_17_17  -7.218785e-01
K1_0_18  L1_0_0  L1_18_18  2.090070e-01
K2_0_18  L2_0_0  L2_18_18  2.090070e-01
K1_0_19  L1_0_0  L1_19_19  7.751308e-01
K2_0_19  L2_0_0  L2_19_19  7.751308e-01
K1_0_20  L1_0_0  L1_20_20  7.273486e-01
K2_0_20  L2_0_0  L2_20_20  7.273486e-01
K1_0_21  L1_0_0  L1_21_21  7.287485e-01
K2_0_21  L2_0_0  L2_21_21  7.287485e-01
K1_0_22  L1_0_0  L1_22_22  7.177172e-01
K2_0_22  L2_0_0  L2_22_22  7.177172e-01
K1_0_23  L1_0_0  L1_23_23  7.216260e-01
K2_0_23  L2_0_0  L2_23_23  7.216260e-01
K1_0_24  L1_0_0  L1_24_24  7.264549e-01
K2_0_24  L2_0_0  L2_24_24  7.264549e-01
K1_0_25  L1_0_0  L1_25_25  7.304515e-01
K2_0_25  L2_0_0  L2_25_25  7.304515e-01
K1_0_26  L1_0_0  L1_26_26  7.211213e-01
K2_0_26  L2_0_0  L2_26_26  7.211213e-01
K1_0_27  L1_0_0  L1_27_27  7.233582e-01
K2_0_27  L2_0_0  L2_27_27  7.233582e-01
K1_0_28  L1_0_0  L1_28_28  7.257783e-01
K2_0_28  L2_0_0  L2_28_28  7.257783e-01
K1_0_29  L1_0_0  L1_29_29  7.227848e-01
K2_0_29  L2_0_0  L2_29_29  7.227848e-01
K1_0_30  L1_0_0  L1_30_30  6.354469e-01
K2_0_30  L2_0_0  L2_30_30  6.354469e-01
K1_0_31  L1_0_0  L1_31_31  6.464784e-01
K2_0_31  L2_0_0  L2_31_31  6.464784e-01
K1_16_17  L1_16_16  L1_17_17  -7.414509e-01
K2_16_17  L2_16_16  L2_17_17  -7.414509e-01
K1_16_18  L1_16_16  L1_18_18  2.427334e-01
K2_16_18  L2_16_16  L2_18_18  2.427334e-01
K1_16_19  L1_16_16  L1_19_19  6.775596e-01
K2_16_19  L2_16_16  L2_19_19  6.775596e-01
K1_16_20  L1_16_16  L1_20_20  7.044962e-01
K2_16_20  L2_16_16  L2_20_20  7.044962e-01
K1_16_21  L1_16_16  L1_21_21  7.633452e-01
K2_16_21  L2_16_16  L2_21_21  7.633452e-01
K1_16_22  L1_16_16  L1_22_22  7.517949e-01
K2_16_22  L2_16_16  L2_22_22  7.517949e-01
K1_16_23  L1_16_16  L1_23_23  7.558873e-01
K2_16_23  L2_16_16  L2_23_23  7.558873e-01
K1_16_24  L1_16_16  L1_24_24  7.609479e-01
K2_16_24  L2_16_16  L2_24_24  7.609479e-01
K1_16_25  L1_16_16  L1_25_25  7.651297e-01
K2_16_25  L2_16_16  L2_25_25  7.651297e-01
K1_16_26  L1_16_16  L1_26_26  7.553637e-01
K2_16_26  L2_16_16  L2_26_26  7.553637e-01
K1_16_27  L1_16_16  L1_27_27  7.576967e-01
K2_16_27  L2_16_16  L2_27_27  7.576967e-01
K1_16_28  L1_16_16  L1_28_28  7.602261e-01
K2_16_28  L2_16_16  L2_28_28  7.602261e-01
K1_16_29  L1_16_16  L1_29_29  7.570900e-01
K2_16_29  L2_16_16  L2_29_29  7.570900e-01
K1_16_30  L1_16_16  L1_30_30  6.318101e-01
K2_16_30  L2_16_16  L2_30_30  6.318101e-01
K1_16_31  L1_16_16  L1_31_31  6.427720e-01
K2_16_31  L2_16_16  L2_31_31  6.427720e-01
K1_17_18  L1_17_17  L1_18_18  1.042691e-01
K2_17_18  L2_17_17  L2_18_18  1.042691e-01
K1_17_19  L1_17_17  L1_19_19  -6.939877e-01
K2_17_19  L2_17_17  L2_19_19  -6.939877e-01
K1_17_20  L1_17_17  L1_20_20  -7.188095e-01
K2_17_20  L2_17_17  L2_20_20  -7.188095e-01
K1_17_21  L1_17_17  L1_21_21  -8.012305e-01
K2_17_21  L2_17_17  L2_21_21  -8.012305e-01
K1_17_22  L1_17_17  L1_22_22  -7.891044e-01
K2_17_22  L2_17_17  L2_22_22  -7.891044e-01
K1_17_23  L1_17_17  L1_23_23  -7.933985e-01
K2_17_23  L2_17_17  L2_23_23  -7.933985e-01
K1_17_24  L1_17_17  L1_24_24  -7.987159e-01
K2_17_24  L2_17_17  L2_24_24  -7.987159e-01
K1_17_25  L1_17_17  L1_25_25  -8.031104e-01
K2_17_25  L2_17_17  L2_25_25  -8.031104e-01
K1_17_26  L1_17_17  L1_26_26  -7.928538e-01
K2_17_26  L2_17_17  L2_26_26  -7.928538e-01
K1_17_27  L1_17_17  L1_27_27  -7.953069e-01
K2_17_27  L2_17_17  L2_27_27  -7.953069e-01
K1_17_28  L1_17_17  L1_28_28  -7.979723e-01
K2_17_28  L2_17_17  L2_28_28  -7.979723e-01
K1_17_29  L1_17_17  L1_29_29  -7.946798e-01
K2_17_29  L2_17_17  L2_29_29  -7.946798e-01
K1_17_30  L1_17_17  L1_30_30  -7.032068e-01
K2_17_30  L2_17_17  L2_30_30  -7.032068e-01
K1_17_31  L1_17_17  L1_31_31  -7.120282e-01
K2_17_31  L2_17_17  L2_31_31  -7.120282e-01
K1_18_19  L1_18_18  L1_19_19  1.967019e-01
K2_18_19  L2_18_18  L2_19_19  1.967019e-01
K1_18_20  L1_18_18  L1_20_20  1.636932e-01
K2_18_20  L2_18_18  L2_20_20  1.636932e-01
K1_18_21  L1_18_18  L1_21_21  4.345176e-01
K2_18_21  L2_18_18  L2_21_21  4.345176e-01
K1_18_22  L1_18_18  L1_22_22  4.269747e-01
K2_18_22  L2_18_18  L2_22_22  4.269747e-01
K1_18_23  L1_18_18  L1_23_23  4.312677e-01
K2_18_23  L2_18_18  L2_23_23  4.312677e-01
K1_18_24  L1_18_18  L1_24_24  4.285970e-01
K2_18_24  L2_18_18  L2_24_24  4.285970e-01
K1_18_25  L1_18_18  L1_25_25  4.308329e-01
K2_18_25  L2_18_18  L2_25_25  4.308329e-01
K1_18_26  L1_18_18  L1_26_26  4.220006e-01
K2_18_26  L2_18_18  L2_26_26  4.220006e-01
K1_18_27  L1_18_18  L1_27_27  4.291495e-01
K2_18_27  L2_18_18  L2_27_27  4.291495e-01
K1_18_28  L1_18_18  L1_28_28  4.263121e-01
K2_18_28  L2_18_18  L2_28_28  4.263121e-01
K1_18_29  L1_18_18  L1_29_29  4.253896e-01
K2_18_29  L2_18_18  L2_29_29  4.253896e-01
K1_18_30  L1_18_18  L1_30_30  6.982515e-02
K2_18_30  L2_18_18  L2_30_30  6.982515e-02
K1_18_31  L1_18_18  L1_31_31  7.638891e-02
K2_18_31  L2_18_18  L2_31_31  7.638891e-02
K1_19_20  L1_19_19  L1_20_20  6.867430e-01
K2_19_20  L2_19_19  L2_20_20  6.867430e-01
K1_19_21  L1_19_19  L1_21_21  6.983552e-01
K2_19_21  L2_19_19  L2_21_21  6.983552e-01
K1_19_22  L1_19_19  L1_22_22  6.877839e-01
K2_19_22  L2_19_19  L2_22_22  6.877839e-01
K1_19_23  L1_19_19  L1_23_23  6.915298e-01
K2_19_23  L2_19_19  L2_23_23  6.915298e-01
K1_19_24  L1_19_19  L1_24_24  6.961571e-01
K2_19_24  L2_19_19  L2_24_24  6.961571e-01
K1_19_25  L1_19_19  L1_25_25  6.999870e-01
K2_19_25  L2_19_19  L2_25_25  6.999870e-01
K1_19_26  L1_19_19  L1_26_26  6.910458e-01
K2_19_26  L2_19_19  L2_26_26  6.910458e-01
K1_19_27  L1_19_19  L1_27_27  6.931896e-01
K2_19_27  L2_19_19  L2_27_27  6.931896e-01
K1_19_28  L1_19_19  L1_28_28  6.955087e-01
K2_19_28  L2_19_19  L2_28_28  6.955087e-01
K1_19_29  L1_19_19  L1_29_29  6.926401e-01
K2_19_29  L2_19_19  L2_29_29  6.926401e-01
K1_19_30  L1_19_19  L1_30_30  6.093427e-01
K2_19_30  L2_19_19  L2_30_30  6.093427e-01
K1_19_31  L1_19_19  L1_31_31  6.199044e-01
K2_19_31  L2_19_19  L2_31_31  6.199044e-01
K1_20_21  L1_20_20  L1_21_21  7.021533e-01
K2_20_21  L2_20_20  L2_21_21  7.021533e-01
K1_20_22  L1_20_20  L1_22_22  6.915261e-01
K2_20_22  L2_20_20  L2_22_22  6.915261e-01
K1_20_23  L1_20_20  L1_23_23  6.952910e-01
K2_20_23  L2_20_20  L2_23_23  6.952910e-01
K1_20_24  L1_20_20  L1_24_24  6.999464e-01
K2_20_24  L2_20_20  L2_24_24  6.999464e-01
K1_20_25  L1_20_20  L1_25_25  7.037962e-01
K2_20_25  L2_20_20  L2_25_25  7.037962e-01
K1_20_26  L1_20_20  L1_26_26  6.948093e-01
K2_20_26  L2_20_20  L2_26_26  6.948093e-01
K1_20_27  L1_20_20  L1_27_27  6.969600e-01
K2_20_27  L2_20_20  L2_27_27  6.969600e-01
K1_20_28  L1_20_20  L1_28_28  6.992920e-01
K2_20_28  L2_20_20  L2_28_28  6.992920e-01
K1_20_29  L1_20_20  L1_29_29  6.964073e-01
K2_20_29  L2_20_20  L2_29_29  6.964073e-01
K1_20_30  L1_20_20  L1_30_30  6.617148e-01
K2_20_30  L2_20_20  L2_30_30  6.617148e-01
K1_20_31  L1_20_20  L1_31_31  6.732869e-01
K2_20_31  L2_20_20  L2_31_31  6.732869e-01
K1_21_22  L1_21_21  L1_22_22  9.211606e-01
K2_21_22  L2_21_21  L2_22_22  9.211606e-01
K1_21_23  L1_21_21  L1_23_23  9.384943e-01
K2_21_23  L2_21_21  L2_23_23  9.384943e-01
K1_21_24  L1_21_21  L1_24_24  9.264348e-01
K2_21_24  L2_21_21  L2_24_24  9.264348e-01
K1_21_25  L1_21_21  L1_25_25  9.339325e-01
K2_21_25  L2_21_21  L2_25_25  9.339325e-01
K1_21_26  L1_21_21  L1_26_26  9.156449e-01
K2_21_26  L2_21_21  L2_26_26  9.156449e-01
K1_21_27  L1_21_21  L1_27_27  9.500722e-01
K2_21_27  L2_21_21  L2_27_27  9.500722e-01
K1_21_28  L1_21_21  L1_28_28  9.259385e-01
K2_21_28  L2_21_21  L2_28_28  9.259385e-01
K1_21_29  L1_21_21  L1_29_29  9.250475e-01
K2_21_29  L2_21_21  L2_29_29  9.250475e-01
K1_21_30  L1_21_21  L1_30_30  6.391451e-01
K2_21_30  L2_21_21  L2_30_30  6.391451e-01
K1_21_31  L1_21_21  L1_31_31  6.501711e-01
K2_21_31  L2_21_21  L2_31_31  6.501711e-01
K1_22_23  L1_22_22  L1_23_23  9.346562e-01
K2_22_23  L2_22_22  L2_23_23  9.346562e-01
K1_22_24  L1_22_22  L1_24_24  9.261994e-01
K2_22_24  L2_22_22  L2_24_24  9.261994e-01
K1_22_25  L1_22_22  L1_25_25  9.254817e-01
K2_22_25  L2_22_22  L2_25_25  9.254817e-01
K1_22_26  L1_22_22  L1_26_26  9.043709e-01
K2_22_26  L2_22_22  L2_26_26  9.043709e-01
K1_22_27  L1_22_22  L1_27_27  9.109971e-01
K2_22_27  L2_22_22  L2_27_27  9.109971e-01
K1_22_28  L1_22_22  L1_28_28  9.103454e-01
K2_22_28  L2_22_22  L2_28_28  9.103454e-01
K1_22_29  L1_22_22  L1_29_29  9.069502e-01
K2_22_29  L2_22_22  L2_29_29  9.069502e-01
K1_22_30  L1_22_22  L1_30_30  6.294723e-01
K2_22_30  L2_22_22  L2_30_30  6.294723e-01
K1_22_31  L1_22_22  L1_31_31  6.403315e-01
K2_22_31  L2_22_22  L2_31_31  6.403315e-01
K1_23_24  L1_23_23  L1_24_24  9.183718e-01
K2_23_24  L2_23_23  L2_24_24  9.183718e-01
K1_23_25  L1_23_23  L1_25_25  9.218788e-01
K2_23_25  L2_23_23  L2_25_25  9.218788e-01
K1_23_26  L1_23_23  L1_26_26  9.039398e-01
K2_23_26  L2_23_23  L2_26_26  9.039398e-01
K1_23_27  L1_23_23  L1_27_27  9.190326e-01
K2_23_27  L2_23_23  L2_27_27  9.190326e-01
K1_23_28  L1_23_23  L1_28_28  9.114172e-01
K2_23_28  L2_23_23  L2_28_28  9.114172e-01
K1_23_29  L1_23_23  L1_29_29  9.088590e-01
K2_23_29  L2_23_23  L2_29_29  9.088590e-01
K1_23_30  L1_23_23  L1_30_30  6.328979e-01
K2_23_30  L2_23_23  L2_30_30  6.328979e-01
K1_23_31  L1_23_23  L1_31_31  6.438163e-01
K2_23_31  L2_23_23  L2_31_31  6.438163e-01
K1_24_25  L1_24_24  L1_25_25  9.523838e-01
K2_24_25  L2_24_24  L2_25_25  9.523838e-01
K1_24_26  L1_24_24  L1_26_26  9.287586e-01
K2_24_26  L2_24_24  L2_26_26  9.287586e-01
K1_24_27  L1_24_24  L1_27_27  9.243136e-01
K2_24_27  L2_24_24  L2_27_27  9.243136e-01
K1_24_28  L1_24_24  L1_28_28  9.308417e-01
K2_24_28  L2_24_24  L2_28_28  9.308417e-01
K1_24_29  L1_24_24  L1_29_29  9.261545e-01
K2_24_29  L2_24_24  L2_29_29  9.261545e-01
K1_24_30  L1_24_24  L1_30_30  6.371398e-01
K2_24_30  L2_24_24  L2_30_30  6.371398e-01
K1_24_31  L1_24_24  L1_31_31  6.481311e-01
K2_24_31  L2_24_24  L2_31_31  6.481311e-01
K1_25_26  L1_25_25  L1_26_26  9.333478e-01
K2_25_26  L2_25_25  L2_26_26  9.333478e-01
K1_25_27  L1_25_25  L1_27_27  9.344408e-01
K2_25_27  L2_25_25  L2_27_27  9.344408e-01
K1_25_28  L1_25_25  L1_28_28  9.412629e-01
K2_25_28  L2_25_25  L2_28_28  9.412629e-01
K1_25_29  L1_25_25  L1_29_29  9.370587e-01
K2_25_29  L2_25_25  L2_29_29  9.370587e-01
K1_25_30  L1_25_25  L1_30_30  6.406441e-01
K2_25_30  L2_25_25  L2_30_30  6.406441e-01
K1_25_31  L1_25_25  L1_31_31  6.516958e-01
K2_25_31  L2_25_25  L2_31_31  6.516958e-01
K1_26_27  L1_26_26  L1_27_27  9.148173e-01
K2_26_27  L2_26_26  L2_27_27  9.148173e-01
K1_26_28  L1_26_26  L1_28_28  9.315181e-01
K2_26_28  L2_26_26  L2_28_28  9.315181e-01
K1_26_29  L1_26_26  L1_29_29  9.218726e-01
K2_26_29  L2_26_26  L2_29_29  9.218726e-01
K1_26_30  L1_26_26  L1_30_30  6.324661e-01
K2_26_30  L2_26_26  L2_30_30  6.324661e-01
K1_26_31  L1_26_26  L1_31_31  6.433767e-01
K2_26_31  L2_26_26  L2_31_31  6.433767e-01
K1_27_28  L1_27_27  L1_28_28  9.277437e-01
K2_27_28  L2_27_27  L2_28_28  9.277437e-01
K1_27_29  L1_27_27  L1_29_29  9.290466e-01
K2_27_29  L2_27_27  L2_29_29  9.290466e-01
K1_27_30  L1_27_27  L1_30_30  6.344193e-01
K2_27_30  L2_27_27  L2_30_30  6.344193e-01
K1_27_31  L1_27_27  L1_31_31  6.453637e-01
K2_27_31  L2_27_27  L2_31_31  6.453637e-01
K1_28_29  L1_28_28  L1_29_29  9.499550e-01
K2_28_29  L2_28_28  L2_29_29  9.499550e-01
K1_28_30  L1_28_28  L1_30_30  6.365447e-01
K2_28_30  L2_28_28  L2_30_30  6.365447e-01
K1_28_31  L1_28_28  L1_31_31  6.475256e-01
K2_28_31  L2_28_28  L2_31_31  6.475256e-01
K1_29_30  L1_29_29  L1_30_30  6.339181e-01
K2_29_30  L2_29_29  L2_30_30  6.339181e-01
K1_29_31  L1_29_29  L1_31_31  6.448538e-01
K2_29_31  L2_29_29  L2_31_31  6.448538e-01
K1_30_31  L1_30_30  L1_31_31  9.550318e-01
K2_30_31  L2_30_30  L2_31_31  9.550318e-01
C_0_1_0_16  U2A5_GND_Group_mid U2A5_V1P0_S0_Group_mid  4.355175e-12
C_0_1_0_17  U2A5_GND_Group_mid Group_602433-081_C2B2_V1P0_S0_2_mid  3.782160e-12
C_0_1_0_18  U2A5_GND_Group_mid Group_602433-081_C3B10_V1P0_S0_2_mid  6.763491e-13
C_0_1_0_19  U2A5_GND_Group_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  4.904355e-12
C_0_1_0_20  U2A5_GND_Group_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  4.198451e-12
C_0_1_0_21  U2A5_GND_Group_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  4.459036e-12
C_0_1_0_22  U2A5_GND_Group_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  4.459084e-12
C_0_1_0_23  U2A5_GND_Group_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  4.459043e-12
C_0_1_0_24  U2A5_GND_Group_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  4.459102e-12
C_0_1_0_25  U2A5_GND_Group_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  4.459151e-12
C_0_1_0_26  U2A5_GND_Group_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  4.459003e-12
C_0_1_0_27  U2A5_GND_Group_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  4.459069e-12
C_0_1_0_28  U2A5_GND_Group_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  4.459054e-12
C_0_1_0_29  U2A5_GND_Group_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  4.459064e-12
C_0_1_0_30  U2A5_GND_Group_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  2.787638e-12
C_0_1_0_31  U2A5_GND_Group_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  2.807007e-12
R_G_0_1_1_16  Group_602433-081_C2B2_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_1_16  Group_602433-081_C2B2_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_1_17  Group_602433-081_C2B2_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_17  Group_602433-081_C2B2_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_18  Group_602433-081_C2B2_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_18  Group_602433-081_C2B2_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_19  Group_602433-081_C2B2_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_19  Group_602433-081_C2B2_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_20  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_20  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_21  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_21  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_22  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_22  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_23  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_23  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_24  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_24  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_25  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_25  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_26  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_26  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_27  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_27  Group_602433-081_C2B2_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_28  Group_602433-081_C2B2_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_28  Group_602433-081_C2B2_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_29  Group_602433-081_C2B2_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_29  Group_602433-081_C2B2_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_30  Group_602433-081_C2B2_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_30  Group_602433-081_C2B2_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_1_31  Group_602433-081_C2B2_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_1_31  Group_602433-081_C2B2_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_16  Group_602433-081_C3B10_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_2_16  Group_602433-081_C3B10_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_2_17  Group_602433-081_C3B10_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_17  Group_602433-081_C3B10_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_18  Group_602433-081_C3B10_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_18  Group_602433-081_C3B10_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_19  Group_602433-081_C3B10_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_19  Group_602433-081_C3B10_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_20  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_20  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_21  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_21  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_22  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_22  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_23  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_23  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_24  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_24  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_25  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_25  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_26  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_26  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_27  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_27  Group_602433-081_C3B10_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_28  Group_602433-081_C3B10_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_28  Group_602433-081_C3B10_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_29  Group_602433-081_C3B10_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_29  Group_602433-081_C3B10_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_30  Group_602433-081_C3B10_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_30  Group_602433-081_C3B10_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_2_31  Group_602433-081_C3B10_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_2_31  Group_602433-081_C3B10_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_16  Group_A36096-108_C3L22_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_3_16  Group_A36096-108_C3L22_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_3_17  Group_A36096-108_C3L22_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_17  Group_A36096-108_C3L22_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_18  Group_A36096-108_C3L22_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_18  Group_A36096-108_C3L22_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_19  Group_A36096-108_C3L22_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_19  Group_A36096-108_C3L22_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_20  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_20  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_21  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_21  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_22  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_22  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_23  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_23  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_24  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_24  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_25  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_25  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_26  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_26  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_27  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_27  Group_A36096-108_C3L22_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_28  Group_A36096-108_C3L22_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_28  Group_A36096-108_C3L22_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_29  Group_A36096-108_C3L22_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_29  Group_A36096-108_C3L22_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_30  Group_A36096-108_C3L22_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_30  Group_A36096-108_C3L22_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_3_31  Group_A36096-108_C3L22_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_3_31  Group_A36096-108_C3L22_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_16  Group_C83410-012_C3L15_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_4_16  Group_C83410-012_C3L15_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_4_17  Group_C83410-012_C3L15_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_17  Group_C83410-012_C3L15_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_18  Group_C83410-012_C3L15_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_18  Group_C83410-012_C3L15_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_19  Group_C83410-012_C3L15_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_19  Group_C83410-012_C3L15_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_20  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_20  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_21  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_21  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_22  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_22  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_23  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_23  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_24  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_24  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_25  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_25  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_26  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_26  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_27  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_27  Group_C83410-012_C3L15_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_28  Group_C83410-012_C3L15_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_28  Group_C83410-012_C3L15_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_29  Group_C83410-012_C3L15_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_29  Group_C83410-012_C3L15_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_30  Group_C83410-012_C3L15_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_30  Group_C83410-012_C3L15_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_4_31  Group_C83410-012_C3L15_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_4_31  Group_C83410-012_C3L15_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_16  Group_C83410-012_C3L17_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_5_16  Group_C83410-012_C3L17_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_5_17  Group_C83410-012_C3L17_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_17  Group_C83410-012_C3L17_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_18  Group_C83410-012_C3L17_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_18  Group_C83410-012_C3L17_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_19  Group_C83410-012_C3L17_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_19  Group_C83410-012_C3L17_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_20  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_20  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_21  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_21  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_22  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_22  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_23  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_23  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_24  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_24  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_25  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_25  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_26  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_26  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_27  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_27  Group_C83410-012_C3L17_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_28  Group_C83410-012_C3L17_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_28  Group_C83410-012_C3L17_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_29  Group_C83410-012_C3L17_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_29  Group_C83410-012_C3L17_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_30  Group_C83410-012_C3L17_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_30  Group_C83410-012_C3L17_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_5_31  Group_C83410-012_C3L17_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_5_31  Group_C83410-012_C3L17_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_16  Group_C83410-012_C3L18_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_6_16  Group_C83410-012_C3L18_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_6_17  Group_C83410-012_C3L18_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_17  Group_C83410-012_C3L18_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_18  Group_C83410-012_C3L18_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_18  Group_C83410-012_C3L18_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_19  Group_C83410-012_C3L18_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_19  Group_C83410-012_C3L18_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_20  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_20  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_21  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_21  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_22  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_22  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_23  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_23  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_24  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_24  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_25  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_25  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_26  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_26  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_27  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_27  Group_C83410-012_C3L18_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_28  Group_C83410-012_C3L18_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_28  Group_C83410-012_C3L18_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_29  Group_C83410-012_C3L18_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_29  Group_C83410-012_C3L18_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_30  Group_C83410-012_C3L18_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_30  Group_C83410-012_C3L18_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_6_31  Group_C83410-012_C3L18_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_6_31  Group_C83410-012_C3L18_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_16  Group_C83410-012_C3L20_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_7_16  Group_C83410-012_C3L20_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_7_17  Group_C83410-012_C3L20_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_17  Group_C83410-012_C3L20_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_18  Group_C83410-012_C3L20_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_18  Group_C83410-012_C3L20_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_19  Group_C83410-012_C3L20_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_19  Group_C83410-012_C3L20_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_20  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_20  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_21  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_21  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_22  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_22  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_23  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_23  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_24  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_24  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_25  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_25  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_26  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_26  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_27  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_27  Group_C83410-012_C3L20_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_28  Group_C83410-012_C3L20_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_28  Group_C83410-012_C3L20_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_29  Group_C83410-012_C3L20_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_29  Group_C83410-012_C3L20_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_30  Group_C83410-012_C3L20_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_30  Group_C83410-012_C3L20_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_7_31  Group_C83410-012_C3L20_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_7_31  Group_C83410-012_C3L20_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_16  Group_C83410-012_C3L24_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_8_16  Group_C83410-012_C3L24_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_8_17  Group_C83410-012_C3L24_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_17  Group_C83410-012_C3L24_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_18  Group_C83410-012_C3L24_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_18  Group_C83410-012_C3L24_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_19  Group_C83410-012_C3L24_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_19  Group_C83410-012_C3L24_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_20  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_20  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_21  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_21  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_22  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_22  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_23  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_23  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_24  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_24  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_25  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_25  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_26  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_26  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_27  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_27  Group_C83410-012_C3L24_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_28  Group_C83410-012_C3L24_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_28  Group_C83410-012_C3L24_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_29  Group_C83410-012_C3L24_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_29  Group_C83410-012_C3L24_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_30  Group_C83410-012_C3L24_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_30  Group_C83410-012_C3L24_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_8_31  Group_C83410-012_C3L24_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_8_31  Group_C83410-012_C3L24_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_16  Group_C83410-012_C3L26_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_9_16  Group_C83410-012_C3L26_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_9_17  Group_C83410-012_C3L26_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_17  Group_C83410-012_C3L26_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_18  Group_C83410-012_C3L26_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_18  Group_C83410-012_C3L26_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_19  Group_C83410-012_C3L26_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_19  Group_C83410-012_C3L26_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_20  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_20  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_21  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_21  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_22  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_22  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_23  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_23  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_24  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_24  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_25  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_25  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_26  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_26  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_27  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_27  Group_C83410-012_C3L26_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_28  Group_C83410-012_C3L26_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_28  Group_C83410-012_C3L26_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_29  Group_C83410-012_C3L26_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_29  Group_C83410-012_C3L26_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_30  Group_C83410-012_C3L26_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_30  Group_C83410-012_C3L26_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_9_31  Group_C83410-012_C3L26_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_9_31  Group_C83410-012_C3L26_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_16  Group_C83410-012_C3L28_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_10_16  Group_C83410-012_C3L28_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_10_17  Group_C83410-012_C3L28_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_17  Group_C83410-012_C3L28_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_18  Group_C83410-012_C3L28_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_18  Group_C83410-012_C3L28_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_19  Group_C83410-012_C3L28_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_19  Group_C83410-012_C3L28_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_20  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_20  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_21  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_21  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_22  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_22  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_23  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_23  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_24  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_24  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_25  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_25  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_26  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_26  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_27  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_27  Group_C83410-012_C3L28_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_28  Group_C83410-012_C3L28_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_28  Group_C83410-012_C3L28_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_29  Group_C83410-012_C3L28_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_29  Group_C83410-012_C3L28_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_30  Group_C83410-012_C3L28_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_30  Group_C83410-012_C3L28_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_10_31  Group_C83410-012_C3L28_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_10_31  Group_C83410-012_C3L28_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_16  Group_C83410-012_C3L29_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_11_16  Group_C83410-012_C3L29_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_11_17  Group_C83410-012_C3L29_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_17  Group_C83410-012_C3L29_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_18  Group_C83410-012_C3L29_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_18  Group_C83410-012_C3L29_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_19  Group_C83410-012_C3L29_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_19  Group_C83410-012_C3L29_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_20  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_20  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_21  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_21  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_22  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_22  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_23  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_23  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_24  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_24  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_25  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_25  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_26  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_26  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_27  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_27  Group_C83410-012_C3L29_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_28  Group_C83410-012_C3L29_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_28  Group_C83410-012_C3L29_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_29  Group_C83410-012_C3L29_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_29  Group_C83410-012_C3L29_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_30  Group_C83410-012_C3L29_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_30  Group_C83410-012_C3L29_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_11_31  Group_C83410-012_C3L29_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_11_31  Group_C83410-012_C3L29_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_16  Group_C97875-001_C3B11_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_12_16  Group_C97875-001_C3B11_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_12_17  Group_C97875-001_C3B11_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_17  Group_C97875-001_C3B11_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_18  Group_C97875-001_C3B11_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_18  Group_C97875-001_C3B11_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_19  Group_C97875-001_C3B11_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_19  Group_C97875-001_C3B11_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_20  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_20  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_21  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_21  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_22  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_22  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_23  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_23  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_24  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_24  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_25  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_25  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_26  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_26  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_27  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_27  Group_C97875-001_C3B11_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_28  Group_C97875-001_C3B11_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_28  Group_C97875-001_C3B11_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_29  Group_C97875-001_C3B11_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_29  Group_C97875-001_C3B11_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_30  Group_C97875-001_C3B11_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_30  Group_C97875-001_C3B11_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_12_31  Group_C97875-001_C3B11_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_12_31  Group_C97875-001_C3B11_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_16  Group_C97875-001_C3B9_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_13_16  Group_C97875-001_C3B9_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_13_17  Group_C97875-001_C3B9_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_17  Group_C97875-001_C3B9_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_18  Group_C97875-001_C3B9_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_18  Group_C97875-001_C3B9_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_19  Group_C97875-001_C3B9_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_19  Group_C97875-001_C3B9_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_20  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_20  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_21  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_21  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_22  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_22  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_23  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_23  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_24  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_24  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_25  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_25  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_26  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_26  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_27  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_27  Group_C97875-001_C3B9_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_28  Group_C97875-001_C3B9_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_28  Group_C97875-001_C3B9_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_29  Group_C97875-001_C3B9_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_29  Group_C97875-001_C3B9_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_30  Group_C97875-001_C3B9_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_30  Group_C97875-001_C3B9_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_13_31  Group_C97875-001_C3B9_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_13_31  Group_C97875-001_C3B9_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_16  Group_E16347-001_C2B12_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_14_16  Group_E16347-001_C2B12_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_14_17  Group_E16347-001_C2B12_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_17  Group_E16347-001_C2B12_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_18  Group_E16347-001_C2B12_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_18  Group_E16347-001_C2B12_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_19  Group_E16347-001_C2B12_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_19  Group_E16347-001_C2B12_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_20  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_20  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_21  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_21  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_22  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_22  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_23  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_23  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_24  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_24  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_25  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_25  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_26  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_26  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_27  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_27  Group_E16347-001_C2B12_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_28  Group_E16347-001_C2B12_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_28  Group_E16347-001_C2B12_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_29  Group_E16347-001_C2B12_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_29  Group_E16347-001_C2B12_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_30  Group_E16347-001_C2B12_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_30  Group_E16347-001_C2B12_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_14_31  Group_E16347-001_C2B12_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_14_31  Group_E16347-001_C2B12_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_16  Group_E16347-001_C3B17_GND_1_mid U2A5_V1P0_S0_Group_mid  1.000000e+09
C_0_1_15_16  Group_E16347-001_C3B17_GND_1_mid U2A5_V1P0_S0_Group_mid  0.000000e+00
R_G_0_1_15_17  Group_E16347-001_C3B17_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_17  Group_E16347-001_C3B17_GND_1_mid Group_602433-081_C2B2_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_18  Group_E16347-001_C3B17_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_18  Group_E16347-001_C3B17_GND_1_mid Group_602433-081_C3B10_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_19  Group_E16347-001_C3B17_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_19  Group_E16347-001_C3B17_GND_1_mid Group_A36096-108_C3L22_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_20  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_20  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L15_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_21  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_21  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L17_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_22  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_22  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L18_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_23  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_23  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L20_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_24  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_24  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L24_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_25  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_25  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L26_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_26  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_26  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L28_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_27  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_27  Group_E16347-001_C3B17_GND_1_mid Group_C83410-012_C3L29_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_28  Group_E16347-001_C3B17_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_28  Group_E16347-001_C3B17_GND_1_mid Group_C97875-001_C3B11_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_29  Group_E16347-001_C3B17_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_29  Group_E16347-001_C3B17_GND_1_mid Group_C97875-001_C3B9_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_30  Group_E16347-001_C3B17_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_30  Group_E16347-001_C3B17_GND_1_mid Group_E16347-001_C2B12_V1P0_S0_2_mid  0.000000e+00
R_G_0_1_15_31  Group_E16347-001_C3B17_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  1.000000e+09
C_0_1_15_31  Group_E16347-001_C3B17_GND_1_mid Group_E16347-001_C3B17_V1P0_S0_2_mid  0.000000e+00
.ends a0002_CPA_Sim_3
