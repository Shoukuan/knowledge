* Path and file = D:\Work\02_SIwave\07_CPA_Flow\A025 PCB RLC Extraction\PCB RLC Extraction.siwaveresults\0002_CPA_Sim_3\0002_CPA_Sim_3_PDN_Channel\0002_CPA_Sim_3_602433-081_C3B10.sp

.subckt a0002_CPA_Sim_3_602433-081_C3B10
+ 1 2
C1 1 2 2.200000e-05
.ends a0002_CPA_Sim_3_602433-081_C3B10
