* Path and file = D:\Work\02_SIwave\07_CPA_Flow\A025 PCB RLC Extraction\PCB RLC Extraction.siwaveresults\0002_CPA_Sim_3\0002_CPA_Sim_3_PDN_Channel\0002_CPA_Sim_3_XW_XW.sp

.subckt a0002_CPA_Sim_3_XW_XW
+ XW_GND_SINK_ XW_V1P0_S0_SINK_
V1 XW_V1P0_S0_SINK_ 0 1.500000e+00
V2 XW_GND_SINK_ 0 0.000000e+00
.ends a0002_CPA_Sim_3_XW_XW
